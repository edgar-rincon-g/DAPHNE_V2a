-- front_end.vhd
-- DAPHNE FPGA AFE front end. Automatic alignment version.
--
-- Jamieson Olsen <jamieson@fnal.gov>

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library unisim;
use unisim.vcomponents.all;

use work.daphne2_package.all;

entity front_end is
port(

    -- AFE interface 5 x 9 = 45 LVDS pairs (7..0 = data, 8 = fclk)

    afe_p: in array_5x9_type;
    afe_n: in array_5x9_type;

    afe_clk_p:  out std_logic; -- copy of 62.5MHz master clock sent to AFEs
    afe_clk_n:  out std_logic;

    -- FPGA interface

    clock:   in  std_logic; -- master clock 62.5MHz
    clock7x: in  std_logic; -- 7 x master clock = 437.5MHz
    sclk200: in  std_logic; -- 200MHz system clock, constant
    reset_clock: in  std_logic; -- sync to clock domain
    reset_sclk200: in std_logic; -- sync to sclk domain
    done:    out std_logic_vector(4 downto 0); -- status of automatic alignment FSM
    warn:    out std_logic_vector(4 downto 0); -- warn of bit errors on the "FCLK" sync pattern
    errcnt:  out array_5x8_type; -- bit error count on the "FCLK" pattern
    fe_trigger: out std_logic; -- self trigger generated by the detection algorithm
    dout:    out array_5x9x14_type -- data synchronized to clock
    
  );
end front_end;

architecture fe_arch of front_end is

    component auto_afe
    port(
        afe_p: in std_logic_vector(8 downto 0);
        afe_n: in std_logic_vector(8 downto 0);
        clock:   in  std_logic;  -- master clock 62.5MHz
        clock7x: in  std_logic;  -- 7 x master clock = 437.5MHz
        reset:   in  std_logic;
        done:    out std_logic;
        warn:    out std_logic;
        errcnt:  out std_logic_vector(7 downto 0);
        dout:    out array_9x14_type
      );
    end component;
    
    component AFE_self_trigger
        Port (
            clk  : in  std_logic;
            rst  : in  std_logic;
            i_data: in array_9x14_type;
            o_data : out array_9x14_type;
            o_trigger : out std_logic_vector(7 downto 0) 
        );
    end component;

    signal clock_out_temp: std_logic;
--    signal data_afe0 : array_9x14_type;
--    signal self_trigger_afe0 : std_logic_vector(7 downto 0);
--    signal data_afe1 : array_9x14_type;
--    signal self_trigger_afe1 : std_logic_vector(7 downto 0);
--    signal data_afe2 : array_9x14_type;
--    signal self_trigger_afe2 : std_logic_vector(7 downto 0);
--    signal data_afe3 : array_9x14_type;
--    signal self_trigger_afe3 : std_logic_vector(7 downto 0);
--    signal data_afe4 : array_9x14_type;
--    signal self_trigger_afe4 : std_logic_vector(7 downto 0);
    signal data_afe : array_5x9x14_type;
    signal self_trigger_afe : array_5x8_type;

begin

    -- this controller is required for calibrating IDELAY elements...

    IDELAYCTRL_inst: IDELAYCTRL
        port map(
            REFCLK => sclk200,
            RST    => reset_sclk200, 
            RDY    => open);

    -- Forward the master clock to the AFEs (via ext clock fanout chip U20)

    ODDR_inst: ODDR 
    generic map( DDR_CLK_EDGE => "OPPOSITE_EDGE" )
    port map(
        Q => clock_out_temp, 
        C => clock,
        CE => '1',
        D1 => '1',
        D2 => '0',
        R  => '0',
        S  => '0');

    OBUFDS_inst: OBUFDS
        generic map(IOSTANDARD=>"LVDS")
        port map(
            I => clock_out_temp,
            O => afe_clk_p,
            OB => afe_clk_n);

    -- make 5 automatic AFE modules

--    gen_afe: for i in 4 downto 0 generate
--        afe_inst: auto_afe
--        port map(
--            afe_p => afe_p(i),
--            afe_n => afe_n(i),
--            clock => clock,
--            clock7x => clock7x,
--            reset => reset_clock,  -- sync to clock, 3 pulses wide
--            done => done(i),
--            warn => warn(i),
--            errcnt => errcnt(i),
--            dout => dout(i)
--        );
--    end generate gen_afe;

  gen_self_trigger: for i in 4 downto 0 generate
    self_trigger_inst: AFE_self_trigger
        Port map(
            clk => clock,
            rst => reset_clock,
            i_data => data_afe(i),
            o_data => dout(i),
            o_trigger =>  self_trigger_afe(i)
        );
        
    end generate gen_self_trigger;
    
  gen_afe: for i in 4 downto 0 generate
    afe_inst: auto_afe
        port map(
            afe_p => afe_p(i),
            afe_n => afe_n(i),
            clock => clock,
            clock7x => clock7x,
            reset => reset_clock,  -- sync to clock, 3 pulses wide
            done => done(i),
            warn => warn(i),
            errcnt => errcnt(i),
            dout => data_afe(i)
        );
           
 end generate gen_afe;

--gen_afe: for i in 4 downto 0 generate
--    AFE0: IF (i=0) generate
--        afe_inst: auto_afe
--        port map(
--            afe_p => afe_p(0),
--            afe_n => afe_n(0),
--            clock => clock,
--            clock7x => clock7x,
--            reset => reset_clock,  -- sync to clock, 3 pulses wide
--            done => done(i),
--            warn => warn(i),
--            errcnt => errcnt(i),
--            dout => data_afe0
--        );
--    end generate AFE0;
        
--    AFE1_4: IF (i>0) generate
--        afe_inst: auto_afe
--        port map(
--            afe_p => afe_p(i),
--            afe_n => afe_n(i),
--            clock => clock,
--            clock7x => clock7x,
--            reset => reset_clock,  -- sync to clock, 3 pulses wide
--            done => done(i),
--            warn => warn(i),
--            errcnt => errcnt(i),
--            dout => dout(i)
--        );
--    end generate AFE1_4;       
-- end generate gen_afe;
    
fe_trigger <= self_trigger_afe(0)(0) or  self_trigger_afe(0)(1) or
                self_trigger_afe(0)(2) or self_trigger_afe(0)(3) or
                self_trigger_afe(0)(4) or self_trigger_afe(0)(5) or
                self_trigger_afe(0)(6) or self_trigger_afe(0)(7) or
                self_trigger_afe(1)(0) or self_trigger_afe(1)(1) or
                self_trigger_afe(1)(2) or self_trigger_afe(1)(3) or
                self_trigger_afe(1)(4) or self_trigger_afe(1)(5) or
                self_trigger_afe(1)(6) or self_trigger_afe(1)(7) or
                self_trigger_afe(2)(0) or self_trigger_afe(2)(1) or
                self_trigger_afe(2)(2) or self_trigger_afe(2)(3) or
                self_trigger_afe(2)(4) or self_trigger_afe(2)(5) or
                self_trigger_afe(2)(6) or self_trigger_afe(2)(7) or
                self_trigger_afe(3)(0) or self_trigger_afe(3)(1) or
                self_trigger_afe(3)(2) or self_trigger_afe(3)(3) or
                self_trigger_afe(3)(4) or self_trigger_afe(3)(5) or
                self_trigger_afe(3)(6) or self_trigger_afe(3)(7) or
                self_trigger_afe(4)(0) or self_trigger_afe(4)(1) or
                self_trigger_afe(4)(2) or self_trigger_afe(4)(3) or
                self_trigger_afe(4)(4) or self_trigger_afe(4)(5) or
                self_trigger_afe(4)(6) or self_trigger_afe(4)(7);

end fe_arch;