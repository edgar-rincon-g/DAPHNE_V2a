`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2.2"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CfYWbKwylvtPqUOzF7uqmK4zs44bz2fdwvpuFLioaHj10Bf6wfz/J6ASNAQkNdzDWKNKpdQVU4js
IClenzy1Gg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CebXybeWb7usVEwvfGGymgkIrvocUle6sj7yT4zEIm4i9uFyh5SaKwhbhgaGQtOTqohXiToS/HWM
ynFvwnrcMSqdNKeH+XTRlujIA0Ur6VKF7Loe/oNp1b7W64pIDqzI77KY5cHbD6/LUNYHhRhvUyrj
A4zdcMalFYRO8xf+eMA=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
u8Q4xIAl+5IQ9LDuPIySUfr+FIAHc3eKWriUMXp2gqpexe2Z62NVfZ6DaIM2aqOTdUbtxTDdWx/r
N6cDE6tB09U4MNuQVpg1LEdmVV/xCvY8plQLPAAGlJJZxN0NeUGrg8UeKgAJM+3UG7oqO3MvPYK2
uEu2XXmKyazbrQFwn4o/Pl1UxWNZ27JWgop7B4FUJ7hnrj4bW0c2rdPL/IA/VeQXe1s0zaCBIFML
iVNxBJimH4+h6uDV33h94bxRWSrwOsTlPLvqFS9IoMeIdYOltcw4WOCF+1NDRRBRSutmgA6w6Zy3
/NwY/HhqUBn4J8PPB+NMAadhztbvmmB+hEXt5w==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Kr3foWuyUzAupd1E7iPi9zkwXkstPmWJWD5y8jxXUVfPbli5ElqScq6V7RUg0ucGB+bMkVy72KkO
4SeTSOOf/ym3a5YrxLjz4hUhYe6QzevP4YGOPnn3xx4PMCtxfeFhvrWf41nqfZI2A5km5njYzbRz
myDkobHiUKDj+k/p33AmOQNwc+nufedrdbd+P43EHF3M5Tu0HUtb6xpzDiK6LJloJr9Vl7k79WzH
7P+G0LKXsGNd+zgC4XU9lyymxVprAjHGqqCpNbmEiI675sEyMbSoCEmrWbLe2OHOjH5/bI/PIZpA
fshbwTarI0jXCu3OniTZDPE2B0OWvGkWYv2A5g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RZ207B06H8GMroXA2sXNxFwurKOqO55VpY16rb2pS4Tr9HrogLWOGcyHRZqG87dS73fhLQ3uQnp/
z+MuAv97WN/bJ2O+8P3Emoh4VuDcKKbOKTmK822UgT5QmUWYQC0fQz3FUiOAqIx2hEnUAlbWPLpS
BxeuGSnBSGSzS7yiWHE=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
asuW5DHy+IbvHkMjfKhvedLnbuvn9AXk03V9JOZXaPKPv81cZQx/d8X1OROFqrUgs4HrYeqmU06t
DVxGtCJmMCxokzose4gcvq9E5GDYqZFvlhpM5eUJDDn5AdhhYyZvhmNBMsl20ooXUX+5XCn2nj2g
LsW5WhaPqAyHMTAb3OgxkQiVZqTcPBmPW4cpxlvy77JMjv8aQ9XKDOAa/gcPswwvZyCr6nIcfUNm
zs1WwDgTP/76Eyyb107vEkjefib52fliAdGzA4pjZTQWV1bDQOIbpAkEsmdgLw3QnCjTwyKlS6US
1/hHaaU13HIvUDEK+pnM+L1ZO2vFR/xwVNuu3w==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
m4lOpjqNlpNhypci9v6ztgXPp8EbVc+wvYWbTc4Da9NqT8uGt0RMFRVdpf7bv/0OZaYMf/f/b6TX
UptCdcrkVZTuVU73QxEFO6D7J/+WcjCg+5/bsvmfi65CxgbzRHQVppl5aLqmLuxW0QU8JkGQEsSN
SQvVG+5kWTqsrkwEoL1Jo+D3UPzb6zU2Fv3NF2nVHp9JypchR5bg2hfGIj9F7cjGBMJqXoiUJopF
YfXjaLc7jl80GwCBLcNqjIoZFqHdR78ckgT2C3YDYcBGy86MwJJq5flQSFUDgbE05HA3FKxzTveL
kdNGVCMqqB0yytu5EnoNcVRZDXhmDen7jTCkQw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OMUi83PSiPalEEiSBiHudEmuQIjQvRZqjQJt6OrYQuPTqxvFanRpm9SDo2z8ueGd6qZK2JiYREEO
5+PJm7Ab8y3F5Ed7H5BR+ZGOwYUlXsWRfV9VhhRymHelQW0bf3UDouo7uViOTsp7ew+BPOjV8hVk
4bYKYiX3d5CUUM/qMF7fyIudHuaiMSPz+1fpIUPH5KiTGmPrvV6HnvyUaB2PIgkE8ddo92BLsQ74
zsy6kx5dbbdBhKuXAlRM4B+x8Vj4+64RiE+kFeAxCPvJ1oW3LDr/GhoGEzyshuaVxjHHtomuL3YT
O2GevzXICki4aNLWfTJJn8gKhdgK4ow4ygRxbQ==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
f4h6vwxLmnvTtsJbdz+fBsfuhR907dusy+EfYSc63f0nY1lD1kEABbKHjGPgxj+4kJxSdJyGjonn
ZbDVMjzFOKen5Q+uU8lnqyzXNUBN9HGiUMLZ2uNK3PPpwv4583hfjeI4VtXw4e/vj3vo12GjSEbS
uTcnLDsCLLfEVhZ8rNECunv/m5BaqTvsQoSDYzzUxVruIEiTLwbt588Y0vxfSpDlvxxYAtPh2aDz
S1TmU9j1pCZGi0jn4tAtRR0Cqk7gZrJbSAFvOkZ8UTl2EFD0U+2rJwSJkhCsECZZQh8X398eMmae
ngTlE3qOYCN7cgGEn9rwWs3pJ1HSHIOJJ2FJiA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 860576)
`protect data_block
TJngYf5PyR1IAgV2BMnW1EqlT3HiHwps+K2tcRwKXQV3B1QpqM0aOZZwS10ZIP79wCc2qUGLL6NN
hIAZKwVpfFTlRm6msimaZvjxO9R8ZWG6SFuy1yb2biDn2xsnL6FtOXP9WADg4OvV6ahesPH+eHd9
HF3+WzX6cGxoHCms6MdUa7AAst64viQhBMjmoA0oq4sGhdDFSE+/bMnJWKD1jRjR6vknPr9vVqao
8TziTnAdmKlUqqvg+BnWsYhKdq52hX6zWDNaX5UCGnFXWkV0aJ9rbD8SMTZpQ1p3QL6RbZgo8PuY
ol4oAOLjoSFpNmybwUHVe/9frQQIqySm6FRzOb9StR05OuksNwWilYhy52UrFYPvbB35P4jFlD7+
t3FIj5HO4XR83dVcYCyAKKfuyik1MNCBR3kHd4aBRH7DGRPxvrLXSeqrcTLv3fYYK7Q95qhxAeHu
YdmjKy0xcohau5ExR5fcupg3YmhbmwHQIFXf3bc7zH8Rs1mPe0oeCwRNfDYGKyB0l9KCHzUvQbv2
9W1NgwAgV6L/b0/g/9sVJlr6x5d2yR4o+83d1Evta7J9uQRd6HUTEFBWvZQuW0cirjC20oZ5zGPN
0Hg4qc486fmEHZRutYrLhM2qi6z1C+gcTfkMhpnwP3kfR8vQaNDLvXuCe9hf6qlidpZMhyssZw84
pImDk+2jsChN5JxT5fcxP+CqTv9Xm8oTwgVR5LBRVvF2mxd9w3YFOi/RJKRCUIMGF6RD1KHR9uy8
tGOwlR9P3Mre0o4bcD9fMgSSQ2khHN5JGJkGZs+ku2K3casKKhQtttGH3zJKrbAZ98s4m12MiLd4
z5yeNOXCfisQGTzavxGKhhkbIUqxyidBGk8hR9fOxiXuHOSnnNID+cTkZIRKjf8TZhHssOpXrJLs
G2nP8KYb9fXkJiF5AIkCO/DLQZPc7+F0FLmH8kkMsKC8tElvYLG4YHMWIn1K/g/GCbOt8kzl80ZS
XAXfmR0GdyLg6cMlbYVlBvDdmEUrigtebpReF8WXVYO6f3AAs0aJCtMTg8c5EJTQ35oG/UHtfdjB
JgqyRqgNku0bGyCTWJ3YvPfFAE/hTxVMwiZdeLva8eDFxGqhH3JHMI6p9UXHE3YPfrB15RMzZ/ev
iL6yHPI5cdJQsOJWN1yIMCigzCaGZkjcAhRIWMv6AfLDurFj0mkhpgb8PpK0hgbkjoWs9CQ4rmer
YYeC+HKYWapkRXK3mZQ4NICA7IvCkKTNAeZ5c0zMZgrEOGkFnySsKkY1V4lDEj6FnMX90AZ+SjuF
t7pGw3JXMy2w10eresgayhd5nfzXhyi2GFE+3xLKg3/fiRloFnn6379TF28MJ39ov4CPYlGkuR5d
WkthkRaf5FVb0r+OgPwStjz8KxgDhL9TrvUHyEKLkI0PBgknwIoJvh7424gXXRhRw0tzUfXC+gvq
+6+O/2KHT/osIv4FHEo5dOA8gut86ISkh+Gp700KpuuiAZjn/I1PAf9y45+j2uKMLal8QhPYjiwx
XyOA2FgmvHSZ17sOm1EDZ3LbOgyYcO8CmWjPA3y1J3h+L5m2+fmoi4PTT8cHpDyVs1C+g2dTIZY3
gVT5ikK8czczGpmOmT6uOJ1iqIaOKoLVeHkwC8ias77EH45sBnDYYBmkztJ9qI4b1u+tUc7uqaJk
Hghnm4rvmSVVHwINTb0Owje4EyfwJ7k/gG3+0ftp2EYbK/Ueq/XJnaQq0GgzibqaEU+kGoauGZXc
Vlic63z7ob9++OpO7XfUJ4KaXxuabEFl9J/vgwRyH+X1UMrKMC/I4BQvf1qrxeKd54ciOHQ3EyWd
h0HDlvi2bbm23hoxcbTSzEhIypDbbV37d7GyEImODlcP9sMKRmKHIzeHAJl4K0WTkEVVN+3JvAut
6IvkisUWwp6CC+1247cAtd6WCT8FZoVQa4C4SkTAf0fxIG97dqAeiRyBR7AgDnUPGNOm4cNG7dq/
iZ7MlJGgUbMllDyLg/TXXFyrpPzGfWwuxJsruK15b3tHbBN4KGrmbmbqpFoHWyug5v705SMsZZ4R
lHnHg1Z2DZcY6o7WKa7+YXrO1OErkx49lRL5tsF6YqzX4oKzgO/RPVOOTD7EiOEBkgSCwFLIb83O
mf3Uglr4ILMNDrndspkuEopoeACdrXTg6hx2GzoGv8E1tngqYcldjPi6MxvX6AAPrwF+1d96YvO6
/O39WJwOWOmy1Q8awt+IHw89qI8TZ2NFFvGPdVgwOB4SXMUl/ztSNz54CpUjT+dHufksvXkEj5wL
wT8HIlozPhMHfKpUqBO3DiIP+MS+CtmEjO8teMuiNvitN+uB76LyTScfaUe99biOJhHle0FK3B26
bFcdc54nl9JQblrbb6OF18+1iTqDL6oCyliASUizPvYPvc/GVyxsBM8sYJVzwyC2dsi9vpi2d2gp
do3koY6jOn1Z6oHRoFMdsB0oqAaI9xGS6vjEL8sx7aPUVBlsJIm+YJ2NZqAA1CMUWIsGUR/ZlwiJ
WLthZCVFY1sYnocjfr4SbAKlrj1k/A6Qpkk/LNxXFcKisYP0Tu45r10kcnMJEiP9u/tXZvBvlUn7
yUDGAvtwUWSCZ+LlsiyQt2l8AWxVHsZCbbk/JX+Qz/m5J8LbzZP7gFyJWLDqRuXJUO9ov4g2upux
vFNuJ8yjHnmERtB+i1/5ccetX2AmbNi2EtgKNxs5yZ4ryW5+DEms61llcbBv2QBIdNM4nGWzdThy
2JmRhcIlj8fpUIgvaEjTid2gpcJJomKJo6TFjsJCujGvrp5jO4opH9/94I+fnUHpF1Ag3veSB49U
726/AtUyGr5lXgCmhXFx96uTixdievtv9XDEaEbPrsSYM8tdUS/zYqLpowqORPoyQLuCDap6mv/h
xZ7+TWu7ONlkgMNljpJcBxd2SgXg3o12GuaN/wseZ8yk1QCw/81c1vc0UENFw9j/oG3SxPGSBnEW
0vdrLU5nDFFTBtfnXzSAov9brrRjvd53DSjsA4CM5GwuAjxdNwU2v7x7VZx5QYPBM+WA8IEjb4/3
fCBug7hhTpSwdaclOXB8wUy+LR52qf++ff4tzpSQXmdjtxHEdhZtX+sCUkwGDK5pNOyARnto3jEW
TrhFVqxex6MwVIwOe1H0Et18Ij4RCG9eZpk7DFhBoR/K22fGhUixxSi49e5aQjj7wa5iTjI0MPKo
5u3jqyuGO7jQ09Rnk4+d06HnKGARYWlpaDS+0ZXcIRSvJMxHqjdI/Jd94RbFgIpP1BMw8VOieAJr
OtJ9xnpsCVE0neCN7/DXW86a8yQWSGhim96rbmUuaRvjPWRRovacX/To1VI8jZ6knJC4MGPu3B+K
T4+rw7LDoKDWpThlKKPaq1WD0DY/GTf9TE14+wP7QaVnzqxVteYoQh9R43ElpI0Ay3hEk9KNirkP
b3jPxCgfRvRC1xaZvgm9WxtBRxwNnGOT+iP3N8K4fIkPGe5YKu2eUhktLU+O9KShT4vQaPbwUtCM
HyJD5XmD9vZ4unRSY4kcrXF7NiyWLg8QNPepxywf8AW7WX1r6Q5LDdiXPIpStn0ndUWsKstx3vGV
czCBoTASJSwmb67H9dabXfHuFGufei7pMdewwvleL/4Qv2Sr2BjOFmjj6gAuKoSfyQErWN9kxJS8
pwFbWWxmWwehlKYSF1aohI4pG7RJ8DTLSVyj/BjD4iU+bFooJ3WBNIN3YEpwXmhMGc1mb2idmZev
bYgJ2vwvDbm/rsfpnmMlhAUzKaWLguFiNqVIKwrOwpNeGcyIcTE+eeuZMgS/gQoSSrELXVRekQvH
wv61taqfPiOzdCDwh7euXZYY26TOmP7rJ2GOAwnXcvfe94/n3oWqDfEpcyvOchV0vdjrYdVXN4uu
7B6W1rKFEshyFUho/y14H8ku5q4B0LUTYpwqbTBo6XkuGNuFY+z2qA5YkSS1zBP+tINWjP5zS4d9
gwI8SW/C7GJ79Kjva4GccBtB+OJrBRUbSDqmnPks6KnGXuDvFMaDNPECclUmurSM9ZIrwlxlufEL
TQkbq5gpVpIOTgY+YoknRv4MDLQDR48jBYO4vUvynEY60jXLwO0RCwlKV9xqIPWKtQWk9Pq4Rj3L
jeYYhi/d0Rb8YRwSB9mUVkzClQcnbDQKNECfen4wnuYVxo/kUw/lk6hLAfBR1Pm8G8+fLdU+uE6x
vE1yfu0I2XDKAZLVPTMuBwCITMl0xVfSJMCs1BwArB8HK9BDypzXxiHtJ6WH0gCnwZbmB0w9I8Kf
Yw2oxvckKhLpgQpDBOEejAJZ17Tzny+6D5u++QamrlBFWP0AOUu7uLW1it5/yiEg9B/G7pVB6wdR
MDJWivqqEicND/QHis4kKHGO0x8dUd6Q/LsokWEbSCu4gt+FLEMB1X/+kxUfIwPEhjd//vpwygXm
UZ1aHco3F2sk153g1gaDAyYQS6sOdYSS8toh67ueC1x2912dY3PTLKAQ8Vsi/kXd8k+DS9jqJDft
yXgrj8ozBNTcxhuNM3tri69iZE8af9+4gB5RMm2Xf3ytL34gFoyNXow+/vpBUrFYXq2aI/eMd1e9
1eMN/XmohNLjDoacX2oxYG6BBe8NqtsKdgRtVQI5PITO649ZGK6Kwi8ijEF9bmX748VfcFeeVuQG
j5HYtd9hhg7sBR44w9eSahpEzHKONpKRRkHRuQR0SqyMgiSdvsJdluvd2qprzafluBKgfS3Bj/6b
IpTjhyJ96GZtwKhSrVuMb/yMyBUNtX7Sq3gEvXbrDLR1TIueM+t/yt/ZaPthmvZDW9TDlva/hqcn
zZni0vaBnrPHl5GGcGXSPiYw/MXff0l8okb3A7YqQ7dU4Y/iI3ReWqWkzQgKdohEg/ggHvJChVzQ
1VKdNRwlEomi+EPgXTjVETjS0jhmdTpZgjHZ+ZH1tMD+gumJLYj+51DiZbrePWIwj22AZhcg7ZnK
01GO5b5/2IKZ3P/6A92X9y9hKQDwp15ZT9dMIjMVbf/tm3lAN/ioh/0riyP8zFtld5roieqYkDkb
rhph4YzOk/5O06fn4QB/yjRxBvOJS8YlZ0ZRcj66X692uwp3lk4ncTX7QjOISTZ0+5i/H+oh0prR
YSNLFKx1DDcWWFHiB8hNAQ0gwXpPICrSOw6q9ftmhWzeR53XrYupsXHf7havXh7WF3cCuSVYKuq+
EljB4fDqBHAmqpVAW1I5lC7p+/eda4npAwhjXVRU3t/8cicsvBiIDUBW4q7oWUFHTe3PBnl0KHD8
iNTF2YKIq/92o1vxxxSPzEBY9poj+dJWb7Wq2B0jI3eRBJox8FEmnjyHILTlnNwenusazRfeKgd8
KGJWd8QBWS7IG4CiMk1D6hywOas6ZrCb9bA1F+IuWSZK+6zquYyqTXtcpzm4rH+TpkVrzM7laq8l
ND6K4UrEvJqGcWaVdW6Ml4a+Jb9Zn808A/vwgWKjjOMmZJn4TCJh0BphJDvDFg8dma36ogF2v5N9
Q6duCwxJSaXN3DQVRotBcgMFLXl94utrIJQP/fUU+if6SrYcd1LCod6r4aMny0m+wAPhEVIzH6nE
Ysg8IZDtbzP+/l6A80D7HwgoLc32N18oQ+L64UMmvYdM4umAjSJtkuCn4nnqiLggSUfqienO5fa8
FRLmyo+++q/u6LUPtsOAxypzZASlgvydKvYJbC+j02685a8KYQ6bnp6cybA/Mq0Wnpv9u+K1cKZ4
N6zmT1yT9fTG38AX1nNHzftG9Ioc7SkgKInrPWvPm5H6R8eIsBx9rFZHeZ+GB40GCDC14ZuxvhPS
wuRU0+I/5yrWGvGy25jROcZN2t9utYCZso4FWzZ5vL+Dvk3Eo7Te63owYZo8dBOOv2l/w9oq0X2d
u+6Un0XDGnzMA7D5ZwJFeXZu6a3y8NDMFhA4d544jefR6/05/atJ5v0K156tCEZnrxWRQ7YY4l9d
+y7WIOfeOhdbwPVhTh8dBmuntl3LcIA02/K6FGhHhUU1vkSPyX+y/7PsHsW83Nka9OG9LEVv3WJ/
rYc/V1HbGWnKG97BaHdgVro/fdXD6W9z74vuLq0GgASPvTg2NQRdhLAM6H0kZ+aPFYS986/CRPXG
ua+pJ2jWUEL1k4qh57Klj47kAYbNsqzysKPA7S8UjO2Yr5y9/swsU8VA+CVICtDx32d6ut/JtiyS
XRTxaoq9/zVVJ+8cBR0s5G1bbTbMLSknl+0oZKwmlOVSQPQbBJ76xU+HgOKIF42IihtAF92Qw8aS
BzklgOvaGJ0lIRYMMgey2bG4/P/svGX6tjnr81IfVRQxsnx8cHneetxXKylbHYvxDAC+D2iEJuPp
PGeX+jhD+GE6W6b8EyGnLONIYoRL3oOjwkq7hW6NgO5NG6+HX4yLadUbswOLzQjAvpi9GmAYOdnC
3+JVHc2RR5cEBTvaHbUvJrRgFhb+4ru+BQgH0QSsKQSQ6pBIEk3psgVGjGYfEEn5RHA3tstfHOSI
/819oXOHlV3J1dQqLXSmLAlgcXrJF910II0opPwuc9/Edg4afSc3EzSwfmOguFflQqG+zbU441Il
CIWbS17Oh90n4fhwVbYDlhi/dqw6oe05vZLBogkN8tNpSp3wPryTiAuJIKUNIXgUmpbbpnvZWVeA
wXcUqeMmhbh6F7dfZTO58oFhwwbrhj4qGrQ7LEquNwUS4qm9wLbQJ8L9sd9oWLyFTgsLDGtoc0RV
iMxMDle8kQSQvWRunRTjYFmll4o4Nt3gBP7JgCIJJjiBziu2+v61tzQOftAZbQY+V3ptV10/5oHf
fcLkYxG45cAx30gAK0Mv1AGihOVQRdnG4awYxWOKNZdS95waAWZB+GDXfQEj82NHrVRgoRI3ds6d
J2zJMQ5xy2tEChmEMk2dlOFS4FNpgmkraOnuWG00vtDx1dGE7x2ViiT+aOYXWdeIscFmwlhU25xs
vvilWmtwyBdyz3Oa2E0wfMuDQXrEhnfQJ1lQpEr+4S3zQ93IOamXkCcpzTXqBBxYzdtxm6nUwlJi
cE/57dp3RPGMcBsAcZQDrZZX0ZGk+XaNX77vE+QErwhKpEuCVbBcjTNccMbZQ6yxcXFzQFJPI0fc
/qqSsrYd1Q72L9eY6VU5z4Pc7bj344lyEhynL0Y2gMfaUpJFUIZ9o69+R+SUltTTO6Z8WJAlPU9U
7HmhLB24/W9tsBt4E7fxZLYB7skRtBp1H2FNDN/x49ZZFdAQbsb8n5v/1jfqCMjv7LJqEu8PwMHF
rdi81cpWs1pX767Mn63TzyTP9QcDtZh9qG7HiaMWnKhHLDgBEub+kMM448r+sgfBmop4kWzkS/if
juIeBmxcqgNe2FOEur5YxftIPLXkXo/m5nPJ2gkVXh4C65kDn9sp5IhtSWrtjqsO2NzrKc2moNyE
vN01rJcgd18LhLRjQkLE55Nvx6Q2svtLCOFoLuH6zXlUXiIF0NPdTLAewJwqd6qe8S9OQUvtPn7Y
3YJ01gvs6/aLAqlAp7/fuc/9pzT8j+HC6Lt6E+VhRNiexPA6BuJLjIAqCrTpTbPccKsRlPj99S4j
ad5wVeid5f8zy8vizJV/tBxzd9YrHm9iYHwTuOvxnbid8qglpmcv+pOb1eJkTqBDUsO5KVgsO+GD
FsqBub/9L+E5r98sd2rpeD/qwSZ9XrqnDUR8YE31Iwo1ARU4mGnG9pHUt3xckRGKYH1F/4JqCXzQ
0TkOxiHfO7TYbD/CXt+R0ZNcjdHjGZziqxIDLP2Dmq7pCmNChKHRl6zrtw3YzRj2AM+3ho877tY6
2p3e/GeLNE9wHoBDxrcyeA0wmAIfVYyoArBEbU9/T7R/453ruAjcs2h78QpRRW9MXbniPbmuj9z9
xTdvyV/PlCzqUAzTsKmEQU+wiiafwdnd9gdIjD0r9GDzDtYk/xP/MCHfJbGkRMm2uKnl2lzG7OgC
CVmGATXz9rPpXFT1owxf9baN5LEn55IFkUhp7cKvW4Ws5Gi3m9Y3wA2CC0cBpZZgTkyvvpWkeGyH
flnortKHZOVKQx0zTlORXwS1cBdegbX6sNPmVzkXPDDZeHWDLQP2YaPZndJnYZi8N3+0fT2iavLQ
ICZwzBVeVKHGtCGQ7rlCZT12RuA7hy7TmqIFEh6RZUNgZ4lsXOT2/idIZWsLAej08sXZp2/xsevV
8khKRutURvlJwI386B2GQhpYZgQxrtpomX7Lv+XEporpESYHu0QWRwStJxcODGnYk+gsusgSaguC
MgmHA7lyK+bAhA9ksQ7KZ5CX1LNI0mpfi6U5BibpLZrGNtdcvSlHLsZIMr1seX3b11Rbr/SeYTcx
5cAGaZa+nFrkJzpFK+nRYjKlnyS/DQAqh1BTRBfvQk0BXeWoPH6VvCG7nVRnmbocpu7mgnHV2RTF
ratuRD1LEwSNFcf+ySPzKUImEcXl56imGtf71buIjOo6AqXiUP8OGIyvoGcXuNsM+o/d4QdKztbx
CFLre180dMI8OnNK+zY9qji8WqJuGaa0U9MIiD2gejcB4+kszRR1c9dVyswaaHpNiUdEdZIyEtoZ
BAF6cJ1ynTjGZv5DQjgBDGNupztesbvQ838oy4CvGv86+2tw+3+QbofNyZ9Wk9KweM09G23GidzG
QfMY7ldOLTKPYuqaPAVFCk9YY9Fhwidj+s/2Foy8kGzhV+ftKX9oVmla7xCzaoV56mOX8fPiZtK3
MJsdXHXv8n8rXbPckHKsvNuIYAw+tUNrvW5Az1eILKXmEw7F3kRjaqLJJ+TSnloFY/jNGfM12DhB
cSF5Wj28bLfeKQuSPQ5hFCAVvuyavGb9LePk5hi9mId++ay9/7cY8ygZJL3u0/P1NJQguCjMXjUG
2wQEhPiJVed05uzktaq1ocr8uoiVyNU/ShR1BXvOAh5+Bdu0MUsW8UdjTs3Q9bkEl+xT1p70QGg5
A/af4IadtxMgIscCcr3P6GlJ5wBLcA99EYid8NM/bUIE/3JxCaVT1i/2IngXldNCYzU3kgjpfKgH
aK7NsQdzuUkQe9zr6wef25jh4vrehdG42j+jBy4BRX3ojtOmVmuV6qNc36cNmujWnWBR1Jv/s3Gw
a9fciIq3ioLb7RT9SjkMifbnwy5N2QkyWR1QcnB9H/KaLNmxQ06dzRNCpN3vBissb7hk5CUhhDfU
Ba1dirRP1tdZBPKRH/djpJcPfp2iYHQUrmKWFF8/n/XksUDI/7J2xQwrGEqqnixghAX1Z2W/8xk/
JRGltY4OeaPRpu+sFe7ryDvXMagiJo5SZxNBY68gzouimpv0Vc5WWHIT5t2RIjrl8myFaUI8Kn15
eBduBEUhVi2dbv8v4YMDhSaUI4OWRX3zg6gNC1hzV71005hTnajWToCd9Hyx5U/EZD+aSSEWozDv
mOmxBjpwKbMml6EOWGt30IRZCF+x++nCaz3TKKy0nTT/mUnal/fTEuFtyXtXJLon83sxoBTJAFgI
WCr++8t9tGnlsugDBVHYhO0kdH1VRda0LeEddgRJja7cx1qtCkbOtrR/5TdhAanPWBtWJwhidHtD
pChDoOU8QOU7i88wU8g5SsQ/X/maxWI1EtViuGPg2BkDJZZOoMXgKa10qo4a5Bjx0lhFeaXZqVp3
azI4kQnEkVQtrDfxwUKAxIjRKqk0eZxKIuE294l2QWp1Z+DTsS0OWb9/61GOdNuJWFgs6Lp9mz9m
GbIqQoNGB4ykCfOINa6OXzKTCrlF5RITeOF/7xaBTNxH/ssguC6J4vE5mHZ7U6YPZARwc5Lqpfhr
IbjJcQZ1soqIOboDIJdtBkcocRsVlFK9WNBPOtXJ/yPqtClMXgyr0i58w5/TvSBdbItvUkMLAOqQ
PBSsUGKw/Yjfr6u76Pk/HCI2w6nnpx0W5WJocOKTxMDwjzm/H1dhwuqUX60dGS2I+hV69iDXPUTE
0dbswIN4tAYbp9rftK+nhXxqBTWUyx4n7b1JLJAU+2T/yMDdtw2LceGDIQWMbxK+/81ovmhv378C
2s5vHNCA1/qtfZjBPp9FrmqiVtwRlZ+oHv+N3Qw+dywAD26zLglCrjHX4Ymhsm2m+ERSlps/lA60
n+0vnM0XDltRtDxT5L/ezP5hPeuJmnjaAAs19V1LPva9t8jowwgA56U1P4p71eXD/siUB2nfdSQP
roO1wW3482Zktg42UyFMKzJc8ul5VFkzc7y75cxEly9tedMe0gcwcaTIgEwELSDIpVW1LmYak3qk
AUdPcq8KXlcsMKL8up5yXVygL7FG4aLZg125YfdZa6BXogat2lk7iEYGnrMHtcqv3Sx9xKrvVVSU
3vwHL//YP1iKHCegjoVpGUeof3gp2uJppttHWnyhsKYHVWwrtmh4rvuRIKNh0x8JMhIUJNtwCVHJ
TKMjfLldmTg1NMxKlCA0lohwhkREUx2Tk/OXXJcIz5UDKS7asFi4omBTgmTR6pgQuDGHbaTYpz5Z
5CZNWc67Qkw3hG7AlVQ4D/39RTBNuUWhKRBgqcPypJx/sb5HuRffSXE0TTedhNnnW7SsiiRHrQDD
fhViH5d3kyxG07fAGlHYGCBTP4GipFbPlaXoScXaGTTEMErmeDXEzU+UohiasRLcwh+cPt/ZGLmT
TFCWSxTbhf7rtJ9t75cI/IE3m/FhqCW1DYNe1EBnyt1C6G084ax5mUrR5CCsH9XO3hvdXucj1mIW
up1/lPJnEhs5N4FO59MGUqEafmPbXeDRuJMj+v6oO87C57M2HCPrgUT66mUckJLFQT4RT5EWihN2
LMv3LqMQCuxrJGdGFeLm8kwTnsWfB52sDBe2DkPM3xojwrCRAjW9HhFAwDWOiQWFxSFOdbHXW0cX
CLF21gTWoCwigELdAPQJCvivjer14KvVHaKxyj7TGUkhaLVmyCYdy3U+4TGgoRHPcqjkUvElHl3g
Cq2E4X7rqN2o7lJRCUyQaTEyYyQ2vo8aZ2agwrsG0KaJdCVVMQTkhDVH0txrPF0yOLN3rNWJv3HF
NwGCXNSSbaxQ89WEYHOXOXkHhC7p3C4/RxTY7rzhxdaEgv9uQ2RhlMuAlF1V6gQ0SHzBgAeOe3G7
0E8bRLpJe/xoUx43YyudxZNxYe6Xp4QN0jXfAn6CpxJkOnyNg6xfIC8ZPhlNzZcc3G2uf0wdFHFj
hbjEF4KUM2nQPeNWtN6zEElD5075GB7CO1crC2/sPoeywdgpIpGX7ocLJfv/tN3ktDRsdPaannM5
NG5idKFgUOOZYtRk3i9EnS5cZTGc0w6Th9jfbqpBQjPXabxFle0uDZz/mORRZJ67k+sIR80mMASh
RkxuDmT1TAv5qIwmaC387GPMEZfyK7wmZsJjZ2oPyce+IXI+c1EzcM+ttLW9ftzLLUCJnbuPLMV7
eanLrKxA2brrBCTim1VfkACCo/uaY/Uws9BqX7OcgJoWXkTCV8q+PtQ4DxlEUvmp5JXZCYRgVGui
Z3j+jG5ApvMzi6EaepkU0Y3WPLcgKOpBUwp/Rvv1kYB8srWHHiYdiXpz3PiQ+Ob1FNSpNBXCKhIr
62WUaAoqALN7xGxrwFo8whMhKFOY2Dsf5/h++vXWN/D0CgHua4G683Q5QJetGCfH6YyvXNRnwaUx
LNfI3Eve0AVsXx8DSwgLjlypUtoSHdecMJVecrEP43RT1FbgzaLWu0y0n49lJ97htlDKhuOOlF/S
riEC81rfSUoEaTSP1vW4ckKmy9qN8rSoijsdGZ2HEXRrlyG5ik2j2Qf0fBYH6O37tX733HgM6mBc
too5QXkoOs8vHXKzQMtD64Jk5YpGtB1IyIOQS0I19zNFSqhHfgSvaUVGVtuuAVu7bU3ari0Ca3+R
zHCWPdwcdSAQMrp2+FU/GT5gbQXVCX1PFPVOsn79zUbx20Y0LR1jgIKsBnIbZ2GS7hu5pMWzhkl0
8ss1pOqKPkEXPjd3fBHq1Jobbzx8OZHb4b9mNker8XKcDn2+ugcdlxYJ5x0uIXSFNr9EwDRbCP91
Sy9119f7Tkb3qUOPPaO8vzIC2Lqq1xa6Wss/xgkasxNm6M37d8Hn5R2pR2fap/bn9obSBlF/tqe+
yzHvi3zeFZM+g86+npbzF6xrV+L1kTs47p4tZRYIrQEQ7dABX/4bvq02TD9BHaNAWttV37aOGCIl
lhefrBYDZWIJXCt9tORgRY1qBZxdA+qWrS5PiXI1OxZCaamUXBGEEfeKCp3lgGsAV4L6chNp2LuD
7OUXdKNudtBNGlMriO1+6HX1pZrzxvYSukUkfyEkHmM0r7ng0CIuRgY58zqCzAZD0ySgUA6AU1tI
nPvW7NLmRlMxeqlVHp/jVZw0N3o4DtZ9DY+rq/+BI5/PVGZhAnq/UrCIt8uP5tG3OsROLrWD/l4R
S+NBLQmZZvRsDsxj4B6MhfxZb5LMMzj1b8+vJHmWH7fWUq/UxWoVhCWV4VJKz49LE/IPtrbtYJcD
yM8+brCkMOTaE2gD9ixWhORQXQfQO+fmVFWtijrj9K6bSErlHIlN6+Cwgdr27ClNIkea6/b6yqtv
c2vrtPBybjmfbC51YzsLWcfXEsdDosP+wV2dA2IwRBwZqadjFPSKpPwJB5s4iET4ml2Tvu36sfkI
7wir+Qws+EZ9AFMckHE8X//PnMJNfDQFdnC9cU9Kff5iJnBtrMvf57qxgeozFLwFeDU6myPzdL9Q
GZFlnc34ySu5YU+KdQ9QVFhWFflCWEFuAUTwN1f1kb2yyA87x3Xx2m+uw919qwWKvOs35W+MosUQ
q5NRFrV63xNhItEJgiErxdirVzbj2yJUINvp7Oub9WTPYyyuLiD+C/HpruJg1noQIKptvT7/rNY8
ZC8ropsjJ4sjleue/xzZAZ9/Ur4DnDwMVvooOtIchmIgdvlPbcGNS1dTXH2Kdm4r8Jkl/Yky2Nhy
h405oR8Y170QE6Q8URdyd0eoRFObjC5o1S+Bu7Cg3ge3ZqKgw5pcXlrf0EiJ8wR4jnXIa/IrlUzs
j7cbXFB9qUagya5rxu6Oqd5B1gB7efqDAj8KKuNcMIB6DaX5alxeQOcTOllcWO3QY9bC75BPpw6W
xqIAEHm3cpxo5XYgC+X0slsV1jMnDhNYfRU85uRvV+9bNONkCagsuF9wWoqovu7CnmR1SEUiD3tH
AiyHGdvyZrIPOrQxXKEH258Y/14v6tWBxZTSmLSNugZg1x0mQMedWwoM5zGGVVL+XPz37AFdD6uC
E9N1FLxS75HurcUVRMh2Vy3pEcAPXG73xGoZ1tGOuP3a+ip1pu59XA3upMjjHsajGPgTFp52aTXZ
IsguVOifw8ghZpvgJyMOiziBkKjjsgTUbrAzAXEXEtdYLCBmMySSaai9bC+P3H0KiEwf8KzCd9wi
+vW6A0g5nS0FJoQHOz8nPgJoFT6FZsRKPv5boH4Xr2g0WEEnr2pFiI6KxBKtSNFE9S1YdAfwsBUd
OU7bgSEdqt6z/FEbwj+lzX3OgAk7ivxPNMrrc3XuWFu4SHtHb+a1m5X5qlqUZAbL6FDEPOcUsGXy
/fJ5uTaI84yj1fKMDlRF1ingH9maY/pXMqWzcudXy1f6sLcgeliQEgIYvoexCKUGFt8kA3vvUxj5
OrL0FAAvBSr5DVfb78m02W0wyUJ3CGQ2MFWbztdvBtBzbS1UwkIhgSbGwvIlitv2WaTa6pV4FTgg
vKXKOvUU+PCYcBJXBVR1yBP/xGOx9il5OiYesZ/4UaqPeLP3UWseiMMRGSWYqXHn0w+vZNP63ITa
Wz5uDmqgz6gcLVSO1isJmr8bjGUHTvqubBqnVSvCMc5i7beUw3tuB6BGczOst1Lcs9JrucCQZf9n
av4cswxGm4IFw32+Jech9KdkXH76yp48xJEy3xX0hWw+f3GuMFIL1vss3Oacp2PGF3e28TVDwPKR
kyrFQO1P0VqQeSfknbiNHX3TRpv2Vq1aKNO8M6dQA7S8sDCx8lu8bclcO1sbmHsZCF0XVP2US8yM
Y+dJHzmTJsQAsi1oyocthinVhMcMkdqtYHeFKayQDuvXHxeSfL+yHfkLW6dcHltfaIXl+7apT9RJ
FCP455xpD4Qn1NlRYXzZRmGfKmdWcJC8arKKm/NvjwxDVHkp6XWsUCFepUrTI7TJqceqkfGtgG3T
Miapj/pnrTBkYaHy1d7deue+35wt5GBtILg8mpPt+4aa3ilO2XNXwWr+VyuMmoqAYLPtJ8ehuvJs
/pXoTdEHZ3TT6MoXfEArwtttuP6KQ/m/BSwGYhHNtwVB7xcDKg7xBOUPPDQ6CsOvEF67RBVqFZkX
ixXHXA4iEAh2n9hMKpI808DOKZzvmImbLgGcbQ5zwmto1Lls+u5g/6Ld0DsylH6BDQ/WsO21CxKE
NB8/8xrik+0ncSwSFWuYb77FaCn6r2SHGVLA+YZ85saLS6THy/sSOqdoZfuxMUQN94ijxTfAK0vN
gMaCUuej4L0Mf4IQvf2vaLreHpIsdPAydNXdY+gIfoF2LVIUKIWzET4JjjNX0Ws0NulhdlpMYets
BrCk88CqyuHmv4XuCKKi+rngHYess8SOuvehQVmfefF2yzrEsq6i0fxIwuHpt+/30XpNrqosr/eS
QdtXwAzrxGmBYpjREU8v1wPwznS0vV9O9O4ajJ4U4UOWl+4ZV0mZv5atexMI+AobnFO94ilCjAEz
0nNQWVyvmVzoodrnUOziGwVQ+W2/u4WhXdpOT2mh/FlGuPLtH0pUfCnQEXndqJ+Va9TT6lisJBG5
WYbI8tOs0X2xSljT0+XAP/umCxAYqxTx5iHSsDzKSlJSzyQIXRfLYKgcTBjYkd5lkMvbb/BEeZR/
kHyqCr8rrjQhhIRCXmj9CL8BtSVHzwRbKJxmNI4T+ndZSrv3tLz28OOz/6BymGFU+T+0ycAi55DI
AYud2ytD29BEHOBvnvEEotQawjwHFOEIBBQAIYGyzeAe+5L1Kk3m276DCLY4xQj6ncdpuFX2CNVL
vCtEh1aWNOgiE7x1glzbe/YOBB2GGEP7vfwa51uGpx39ztTtQUz9LGYJ/Q2/5H7QT27RJ4AVWAnn
yrF4MXaUJk53YdlzG36dcXb48zRXGVdiWFAAOzBYVdDM+dLE63lf9n07mNmuAgyglOxiNIrXnRD4
H+TI/BVdro4nbkWyV/FXnLeEYtKbEm5ukktr43uyTEOSLLqymNSrOn9DUOmLaDVp0wLv0/MgRfMc
4ZGMxvCI4UA2gmNgPdvgv/bTDVBC1Bx6/IcJYh5aLD7unP7AzXFi1+QAGnrRyDgmhrWKOt9fDsKz
Tj98UTU1FB1ekBULlTv1VWC1Pxuu3CGjGHlqrvpOXZcI/99uKB4P4WCQI+ZvpApRqY+V9xUC9sLD
wULaFqOJmh+0ks8x6K/aRhHBbhajJu+LrqoZDiBtSI/W/lQw+Sy+aCS8LkRkFCkTmxxMjN4YIXn6
G1aOEvMi5PCDkhBlXMPPQSwp83UeDUVwSZUrrosAjNeQ59JX5MFjAzM0V1u5j6AFQfVE1lkTrPUE
notaH1Vd+fDZn3H5rO05VSLuUHxoz+HvPhZd3jbntr8cyxODkbkQiBwleWowvUvz+MlN3Wok8+tY
GVxD7cZCNbk5h6vvD4PxtIOdB7TSjoJL6NPgLL1dgdNJaqrRDsDmobYzLcIsnomwXfbyC+SYdSmM
Knt2BIjAcejP40ufbJ0XTvb16oll87w8l3iJcb3uTuEo8heQElR72g8brqZE7o4S7AUdurDlBBfB
K8izOgOJ70SrDKd2zlwZDlyJhcSIVXOtdKZ+g3oKReh/IhWS/4oEQK9ALMZBeB4zZZ9YS9tmHu5/
bouiS4Zd4eIoKa9GiCVAVjTYy8+hEpnWfccFmMnMkrKs85IwdN/NJCJHFj3Y66g+ij3qiL28JNRT
9qDwfUVEYELtM85HyCGhEZ/GozDCqiSQTX2oQKx36psLBQCEL4VYyRCu2zdsubz9VKkJweow94ZF
0vTXQejCWbJrVmy5muhyNqWODeOXOKA2+OtVkfnS/zb4VuOelh70fwavawmXGB+sHm+Dbd8sl19k
q7A7Pqkwj77fx3lE+0FjtwHWxxDtcxnLX7gzd4QF220m7METd9BnoCxmxLZvIYifv7mr0vNOzCW1
ujAn2nNMXM50A6hBq7l0PqXB8aKM54jIktjAWX2x1KFExDqhh2qaJx3tYmqYe3hpeYmPZJLfIhb5
lMolCPF78a3MbSucUNAB1bQuWcomfHBR8+HsqXUiuhB3JCnucAVwQHizBZLYcsbjprI9ya+V/Gr2
AV6lyPYFCMXV9lK9X2c8kh++vga/Q/1eVNgZm3bwMM9BZ8QwbugZASVz0vNdGAn4h5CxD38l7s81
Yv8xOLF3rIMku7XVuVRFvLFD6QkIFpTTI/lIpGg91WHe83xSd+J70N5YBeEgQ7dfikeEPqaZ6fH7
EBgQw19S5E17xdQX2nScxKrV+MV9foYeLsx7okFe4eis7AuvHRY4iiinDRFKNBk+8U1hrx6IM1N1
9hHcJ5Los7ikW4Zlvkv7XuPPojIKDCv3bHT3qgKOW3UsiVKwu0hCM0h0Y/bSjSa4UN7Cl0vEpdBB
FZ09WnlRiSezN7XKVrVc7n4713x/iIofx37ROvS18Txv5u1pfJFRxx1dwhYr6EK1aEIHw4y8jc4M
SkefSV9jZNqHlAtpxd0YmI7dHxkjinlIUAYT1n58jgOiODmsj5L0n6B7vTWGWkAu+fwZ6r+0CH42
y2Ou1tqBrKsHv6508LG2NubLmsu5i1RDdGm26vcZt98K74hBFkmQNONQLQ7+znk1eDRvoRsbnhvS
I/Pru2jpuMGI6M+x1QTJsIJZfSo3+uYQHCvI8SmjCyyW3HZ5VeEQYz50VzXYZZh0KeSSWvR/UPbF
NOULClVUKNStFss4/zYahY4ihR92PeeaAReZvDBrWIL7KvOE8WhaNVu7jBOi3GN7U54miV9jHLKZ
pUe/OiQrbl2wmofCdgTV4JfwCiHE7J3a6uOKphE7cUIUtlOvfgDirA4P8c9vU3utluobTiSW/ub8
Xg83uUdgKO1lAYbAcLFyJoTFYCNw3ItGYnZz8JxOjfHHxwUZqEIAyKj4SvhwuK6b1svlOrFV0sS2
AQaOUhwWVmNSUz6jvNYDwenqhVLYH0DjixEnvO6YUlHM2f5EPaS1qPTzn2Ck1KiwYX9ceg/ZmgeD
lfEEsBWWFVT5ae7eGi8W5Q8tcANR7m+ImeVm9GacCEcFkl0P6iOUCssEARxtrNDP5CioQwdgWGim
YIbT7N8Roj9UY1opcs0uP49v256iiTG8PiIBKOo+O99n/SmLjcUjGWIqIwd8Z/ZWuMSfWaiOw944
a94iL9Muq8tAOzQIGTN1dDuP5GUoXJXczaP/GrwBTN4M+Vzty9dNcFvRYAHGkzn+09uCYKGvD+vZ
5DhyxDvMFw0KuoqAu2VCxtPMU1Z2pCqbaI5x9hk2ges4y+012YxjDzICwy9tWQwzNrmK12Y4xIjh
zanJ9JD02cd9Q9qkbXRx898JKwfMw502RzpeIcq1TCTg2ZZqif1ZSELMn5Vni/QTfpxtevZxC9Gr
dmAabBpp7NLW4DzypQBY50FI9FaxJItSJShqkJd6iG86V/FeVUww5mt4GPksn5ew1p8J4a4Bvkmj
U17EEJ/TuQy2PKuu0UvibYBcAicQA/nNmgnoIa1zuWj8AwGRnvQxh0a7a2/+YKuTvVtELjyZN/No
2ODRqn6zNiODsF2dFjXYwAolr84/D+gq75OxGhQ7P+j5YK51DGn2fiDuzr6wkWqOGAnEjf936HFp
Qreh7aZBZfl9eEl0MynGEScABDm+ImYx7MdMPwzYd5rEmtpb/2x+U6ChIlOtG9WDvvYDcv+9IGAY
pYbFnEVl7lZQcY4wUh22fYLDIa9aTFVykvtImXoqMJ+inBvLl0DImttmQUobmcYlNLedP0HNrLFB
29vk96sj3dG4r7Mk+A7pjzbL80//a5ZxCD3/o2o2hlbJW6RrEB1SEVBWvJ1NqlfYGW5sHXszlnEZ
kSf/wSuO2sXQLIMlpWpOZZN+fZXGQZbp4774K3LmeiGXOCp4vzDxmzTz7GemHKlSjrDHUYeKG1rp
K6qnkoOpc+d4ytUbB8bf5EyqHMSeeoh5oi6+sH7OkT7LRF5yFwgZWoHIXxoWhwEGYt6F5hmv6pbH
3WYrXsvVkUH/OgJ98oKf/o1FKx+P/M2nqAFMwouVAmSag+mjtCDhMu7eQVT/mvHxqTADf5USk5bu
SQLa9spQshUpMf9bhcysUn094F90S6lBO/iwNMpHKCv+YILe7mBcaos0IAg+EjYFBqqWiEBqvL5y
KbBm7TMgz9OM7kLCToIwvHLVUQjsMc58V7iNKzGL0fYAJ8zWg42vPJyv+/skoScfVWMorLCNiBVY
PXKMjfshyMzsueGJhSU/KHtZxFxhpB7xlFEsw3SffqpY0Y8KvNMLKqyFDis82UgIHGIsksmxWG6A
QZYddGBTO5LbNkbxbA075otkGhyP8qntklC/aEtZzLnyuJZKLeJt9bPbTEBJQXnNKtwW1ojl81Bt
z0S3b76h56PB0VhoBzZ6RZ/+3w+jcDr/3nfKkVA1GbmpEXpbmnlA8KtSMpOo86ccqAPK13k0E9cb
apKu8S6cZOVtCOsnN3hY55NYuV8CLqCyhV2ZB1b9Dkct2ToJCTsg2rxdCKJNkc60ew9e26I/w2CU
OYu17cZkM363Vay8QcEezrHLrYMnJ9WUr4VArpt0/E3LwtbwUGiF8217breZddHxhJahxfyTDakx
hrh6xUm8O+Bp3kotSBvp7x2jnjRUnb5RZ+LZOm5G2nJ9ccQ5eagBzyJ/wmA7UFbj/WctOKheILzq
Qo7DRl4gyMKNkRQHXC4LjzzPg84XbSW9vQjmS98vZyr9HqFeru/NY6uGXOua61V7WHSd5WsQIWKG
WU6iJvrj3oHdElHq4Nem4+Nn7dlrHBy6bGEOwVvfKmzjAPixk2Op1jk4qS7+mtqpqEA0EvffIRga
AZbUXdel9/AjdQGb8pTYVBSPX0ouh9S8funeEzdhPkxprOm0mk4cSA3DU5r//HM7BeX2jqaDrGKZ
A0zmj1thmIrz5B7glknC4pDgCJzhWgBJz1p9uKmYJKsyA1FxXCErsld/u5aW4e3Nir50EeGm10D6
/TAARt6CpFv4sdUwIQN0gIvVnSKV8otJYlfiOms20n4RKNgiTo9ytSeqYTZaW+oYUTVToRqTR156
JYKmSM/N4vdbJWT/aqg3zax5LJvJ0ad2hk4nJcje0ZRUGBxAASb4B7/qPI1T1W3F0H7FDIcuB5U1
eeTScO1LA5UXbG9JEYhulj+cl9/QfyHjXwQsfdHlWf1Gc32ilpMB5QLtFMj3b8zWNA2pLCARmffW
OKU21PxcGQImwAMPrYQBJ6BHzz9jLcD4GH37fo3WTuVm5gasJl9jIr+YSqnYxU9jtclyZ/0NJ2Mc
r6Aeaj0M/dUuLQbSNzrrUeGeK4CP5/uSbYFGeX15oplLKs/YwkXqtm3Nyd987+41AEj1ZaC8cKbc
QS8FWPYOg6qU0Wofq5DUmAWnhYeoUz233yi0gjCZ3May7dItRhrXxl3k1h7vr6RA0djPhmSueLQr
pwmBbJrfBWsIRyAVzcNl908/PxtwEmcEKpFVw8IMGDANVYgjK0MIM/qT1g2rR/tb1RJPtBRcxFfW
7cJU+yDu1I944XXLWMRteKVieyyX5p+9qlwn/HX/zaOkDa1uXbsp7xek1yRvNLng/75xMe53fOTD
3X+hIELcHVzSiUCUJpQetvMazKppsLmZjst8oO5b0zQbZfvgDJ1GrWyVOAFYBX7mlJSAYqJI9ix9
bnhoQzqZgvjmIMdm005r5iEQb7SNwtF8DnVjX5Ln4lcJRV8AzWJoWY180w9uvB3FUBMMMmh8lnM+
e43qHhxpzZwrzQBYR8PzJ22DbnMvtSd1b5Lw8MMjyz6oqR2kbXI65HXZ3rrdNrg13idfWuSa2o9J
WzQOeiWb2Ewib97WicoADtq8BIRHXgiI++S2oqLqSK6FeT0hCWLrwokYjnsXRLVEY1x0TpEdiXuL
7ESRWihO4kdSTZcdsZfIURtnNAljQML/3sn1jfKkt4lxLZdCW4QQz2TaUw+XYoULZeleTzWF86TO
fuUuNuQix0jfu/KggL3+0YWBVi9FfYywURe7+76EB+h26V3nF4tLZPpsA3IjStOlUI4c53SJblbN
C5uSalCHK2WeENmJxTCf49dvg1DxewsKe1Mx9EJXV1K3y2qojpNQHy+V6JenVYghLGMk18oVIT5Q
TqBOKH1l635vYf5LUHeur8Ve0rlgKCH2KMg0hocVkr6qMb4J/x0jGhroQRzGSW+dJbmXi4tb8OKV
y0dHBQc9SeGqYrSR4uYAH9VqZQqdpkAndjJUTD4XCpv41B1ery7bFq7Z5nvOH3Omtdb8sB+FeOAi
6eov0R+6xcT8JfvLXJpQp8B4jxnsJM8ARYaBSny+QVNCuokhwGbOurroPx/iR0cPNazWjf2vbWtI
BSb6IzLxVSDO0ydgAfPx6RwzinlsmUwFaICBrPdQ53mWNf3wQLvbUbFwsm4LtDzGFoTOscF4DEPL
9gN69XrPHc2QJEy67ZrQItyQlDGQaV2D/RUso/hCl4jW7n02+bDwU7t2O778cRBz0+pA3PGvOo6O
cJB1x3qYrvX3GIbu819Aa/9PSgqXA3zn+wxBEBfgnzmgmkX07k5bXqu8y9mp74qEtYxLh/IlSM+F
7kwYz+ludhhCRCs67iVLLuydCOm5fBCqg9EupJLzOcRRzubdqRSfqvia+Zjlqx0f7Z4JkLsu5CB4
rEuaKRvhbZPCRT1kobCgdq6UG4GKYz8pkW5Tuv9xuzVNPDZ1dpHy+32glaUAm5iynPWdlVocozmE
E+rJ36By8eCGSbgzVq3DwJ7p6KSCagiKxrEZf5pV4Z9hV3MT168WE1fVZxiWq4vr6xznXNG/1ONL
BrvM2yds0QIEsEVwVxGijYyT2h1iCn5kP4wut1WFgUNFaALwNyZ0J3sBfiyer600+jeVAesPEZJa
6sLW+LPnlOe8+JKUln2kVTE+qrzfPAmQgTEX/YmjstITNbYdSzJJa8n293wnF405IEqIuXcJBFaS
GYTIbzEyW3GbQt/VwQeVijpvhmPrFhVv2OCks1sOevFaOAeTHlLekROqGHfHPpTEYrdJKGAvnIKw
1cr5+ub0cgKxNkt9i7qJfY2VPQ8Jg2xnIZpp1bnbY7Hf/g8Z7cWyb8m9TxbY3ItKeu4+nINJWk7f
u4IJzHXbp68bDSMR0nHMMHm/QIFuod4Hdv8aAAx75VEbL/NHMwD99qRkmrX6OpQNOO0UdRsU1eZn
j4YQTHaIVYlXW0wzTLioicyn9gIhiCtlWs3ZysISH6Hqib2lelDY7U4YwXJVJJpKELQ3OVu1uroE
EzvLZCU+E9AbcLJFvQ3kDln5+IR5lOFY/2P9i5Sx7TA2rENBF1Z6fnfGY7wLxnPe3Klq0mmgG7E9
gH37LfkYS/1O2mZfoz4xzsHqv+dijye68rZPpRJxsp2tKhQBKiChGRE1M5Rk5tH+pFtRgTaHhWxu
Wx1czGv5NBpVBvT7FWs1NGEQEg2yQ3Yp0vgH/kGrAw/8pEm7b0WKJ4yJjtbS9TnsVUOWlQD646S5
pH0aHnbGCbuAY4+6pECzPMk2QIJxe06CXoqRsco/Sn24F1osnogHkBjKiz3zfH1fMDgugg/cXJ35
fzZkOLJghe8pzmfeeqCkUR9StMvRU9WbVxfr5k/Ri7QiT8F6DhQwtZOa+tN7WSHRM5rXNFt/hBXp
u+o9D/wvKyqFzHlDTPMXzBgetPn15CiI6xzg6cppaXgaYmuy3CyHURVsFAn3IhOwwgnAq7mIXOYp
nLrGEWA8YYEnFC3ldTv3VRx3IBVZkFRazfWIlITZESf0Mc0KN7mxW2YoMKds+8xMqTOWsLtRtMjV
0e9YWfiosxVZ8xL65uj+0pZXWvNGFxk1vw9eZh0adH2yvP75r+VRmfiQQ0UiKiwUklYneNU7mdZF
AY7YdKqdG4QXEQq3/Wcag+Qd8DfTt78Cp+z1RMtiIoQVpzlMc+12NHNACWPtLInJWMfa7b+qPBql
RjztRHGNsW9apqP04Sj8fAQqT3suuzAKkFvxAszQtyNj+myneTCgWqG2KLwsVCtSFhOfogc+w40y
U7ZMVqNNoR1hv1bzN0DK5nr1tMda2Rs+Xx0vH211QNCf1EcK0EKfs5vSHqXCWCjBgBqXD4u6/FSk
Vq/y1ke53pAfgNanHL+XA2UVV/nf9U6R3vrYnnNw3ObYSQwFE0SpGtpAV1OZb0Wownv7rhmZmPog
dNFKD8yy1aPOY9cYcKAgXF2aFdZKkxJ31QGjbrMOIbcuPQV88DuwDDzJFBw+sojjVFWaBvR1ezJ7
24RJWLv2UXDx8/vX/j712lvxNFUEZIg3dLFzAymvyOU0ZbG+Zfrhw03XBi5ks84lMsCNxfueDh2R
PZs+d1UVdz7qmOM6K8xBOakGaIcDwgerLmpI6Z7tcHUNDP1FvPiRLMiCLUQ7EWxfk5Rl5eOAOPZ1
2FryVQjgpjqfsMBlBdIP1s+n2U+lRaXM2kHvLUqT0w8kSeM5WNazZA/zcJIY9cE/ILnyLKp1S+FH
sHVp2a5bmNkGzm+BrdbtW9cMQj9mtIQSJJH2LK75yrXtwXVmp75j92rxkHlqgiZle1M+Ae0f8ZXU
Pl2m30f5W3LrXwzzNPhLbguSESyjmenTR+zLX7feLB2KYWzmK8+Ib/Wry2/eZqa2DiRt+ysJs2sp
zHwOEepJ0a5V7One+PE7IVwW28ahvDo+Z9zvd/i+tiKEnv8zvmX2sJK0AXHr9AN7odMxScsQ1bjg
3M5MQv1DDiOctO7oCYjoBqJ2CcdY4tt+jbQfHGzRmMSxe9xD93e1m/KqSTTvfZYQwTq5bJEw0u3i
n9iMy/AVwhziNpx44k/+oyRL5DTki7FmTmyY4wi/gHeGkCjxJIGukd8S3EOWy/E506H+fI1eQKM9
RMWpHSFh7dCoOkFP+oW9S+3zDBLdVHqlX5aKjMAe9I9CGJTN9M4h/toM/4kGzSa7dx7HMOptH+Wr
NqO4byLiINMOAZBL9beCp93iyckFnqZViWigfIDKrVvXp9ngiDWvCjygXCpEI5T9mI8WkVbOVmHW
rIYtkxs8nRbzNOTcSGsGyNc1pLpNlpPhNuywxSukAUc+s23cC8by8LYryA2XPe0j8/GvXR4yFEht
ZaC1gs8qRNI7dAwGJjvVcCqvYO1cZ4OHGvMI/ckRRy+LUQ9ZUrYnlyzU1gOOjR4dPMv+6d/dDy7E
2/2gfUF/dOsjSDCpu1keLgNOe/UgUSqkjeL6t/epV7dy+NW5NoRcu0zZBnclT8AuZE8nLKr2Tp9F
oNIVoYMkpM/pF62yzgyf1h8fId9+O6Sodf46BcJwGS3RC1HiEjO3wIlUgYCPD1uc1PLMhe52KOSR
kGjAFbzgldBjZ97Ii/pq8PQJUfwn4gxtz8rUFo17ZoZuZaB25uN4pJiWtWI/iHJdvEGZodD2F3QT
9Sq0PyaNrfehgnyLKV/VuhHEugbNtGvur+jAnnUaHzph0BnlGsyQaRhihzdVPXq/dnEbhPcsLlC3
DUkexqfrxUSCw4fQ0VLAbbWTicaN7shKdxRHnpbYmRNgBv3127R8Ui0tkZM5X5xal2Ujnisg/dU7
h3Pw9NouYIjeq2DERjABaeX8N8awMC3gWKxdjUpUuul8z3ekuS3ac6eLmSkP1yfWhmaD/bOpZKjw
JtQGVGEJWb35E84f6YqLG313ihk3k8LExXbhRhv8DZj3xSN+qMxqfWp9jKNyE1DLtw3CXITM8Nzq
GMrqGEDZyAkkuxU8T+UEA0fSwcYcIlFmPimDlzV6PW7JBIKqAUcY+ikWIJd8sxvyL6ehmxIhc0Ew
dIvpAf/tQmyLqZmyyBbddQ/KbhZybHtsiQpXAXHmT0mawScHOSI5bs1z+IaEnYdxKSFzxLIWEKYF
GEuIBZRJAdGnWeZmKaLPARzwAfCHazlKDauyKWuCwXxSZtrWy5eKT2s/L0/bXgg7WRArI2EpvFlB
Kk0+3MJQVjvVxo0iRDSNgNDBQKK/15JFozeuX28XbJHfrC8lB/OG4ni3M8s7YwM0v2Uue2H4+DkH
PzKZf5hIt3Mzjriczmr0MjDXRrcKtwE/Dg9uIOMgi0PpYL0JVtAigzd/e+TuNLLKhsc3r59jKADy
9SteJTcEf3E4uVlJAj7AF1O1nPlJBgZx6MpJ3+eypNeKbtPQtSWgemKyx6SKhmgbsB0RC4GuAF5b
PFp+t3A0GB/C6lskaE8X8wIyL+/51LpfzTGtJwNLrlSITLgBjQ8n2If148xaqDGY+mL5DWV46Cxu
30Au3JTjuBFamsyfoRtyYwxJ8dNa6O4NtiOe9diClmpETTvUKK0cf/w5us7d8JtU4/Jnt+pC7TAw
LpRKJFbY5rRPOuKfDJ7RswMMZPRcgcYAUG5hrKXHT5tx6Kod+2mZK87OZAACqZ3mmFQUZ26qNoHC
Cx2FFa8IcnNsEa3SwPH/NIJXzoZGW7dPAfuEXgkzFBr0EWOpwuQ8m+z4MumONV/m+IYCg3Y1mfLa
9COBvSZIidhRywzi2pBGA/OKjYrS8b5WEixCcYbtHQ88JrqP4tVpW88aUejiT2UY5BGdaNdnSxGR
VOfXxHd6gVgjFojsmvb2+/Ze48Nwuw4JLp4e4lXuRqbrdb80zp18XndXefS1uMZ/vyzyRhXXA2o0
R16m090qJCDO7HplV5CzmzG6B5gqZ0as6EaGBf+t1crOLS6ZXiah9erBA/bN8dyyF5iCn2quRmp8
4jTNF/IGJK/AnyhzUzmqNWPk9bGZIbnRh2qBAQXHPAyXIqBGSlKVeil0mL2xpgL8lwA3dzs/CXVn
4B6sqSSI0bPoIH4N+1L7SOJ8SZkjexjviBP7P8jVOMLbYiAKV6H9l+FGgNRK3/KiIutJB+OOiHMN
vOxgx9WY3KSBEjdgvUxioyR1Gca8QXf2nF+w/r+Nfp6bJgWpb7SMoKSERKCIz76E01QJuiZ9p64/
zcS64Slx0GmrRj1zUa8dUhNSFlnmmwaSzAIE2cipuQ+87mgMsDJi60KKzP6SOThLKhb5kark2Odk
RdoCAm7Q8Fx/ASM1fzrQI+n8YKVmFRi4j4Aa3L27tXdu5Udw7QnrnRhe7l/6JP0T/TjJAfOIBWM/
7Igwk/fTTIYa0whYjn+R3/LJXOayjupGkLR1f5mHl9daKGBJecnGlPiJMyHpnnJwH8A1dzyrAeFt
3zhNHtuJT4TtsyF4yRDVN/JvpVlxLJDParX09+QPgHmvFPSXPr6CVBL7MTkqGStWFyq5W2AC96OG
+x+qTfrR0xncgWCthICSFUPpB8HBM7z9wY8jAp1CjdU5I3AS28BpOXdqedVf6DIuuiNSiwYmLhxx
bC+DuiJTsYrR6uOf4vU+fPToKhe4jAKCFJPK4P0Y3xPcrHrtE+VXkeQ0NUK1jYVgCTKdp2nNaAXx
5vcBORDo8LwoxXk13YjHF1pxCEHWH4EO2lqAqSZfgBBfKMU1dwP5Ox3b6ybkvSfluhzmbgKEFBPI
q9QkkfLS9W/wiYVahizpr7SEyVdJBlcazgrPfYsIoqck1X6fNKh1fra0l8v1dO5dumxIlj9MJeKf
p2ypi+UQiZzwG68Wwe7HV//wW4f/WSV9asJPeNPTRjK5VcmHVADKmWs+GAXXIBqst8bx6ipdgNeq
nzPwUT5ScxnpKLw4wNchs280tC3v8A1GAlONWHZw7A/eaiv8s0G9Mo9LsKu+O1ZiLaSEHOfC8Jla
mBwXLtx//hLD5ZBElzi0aWPsuo93kuov8Y1P0Yo+Oh4OLVB2g/dk+d69MGEkzj+jAZtIncZpuKG8
Z++uIbrIQGV1rTntQDmPySydYBSlph6SgAKWVIzIyz/h7gKQ6/gfNRWhrXENAnWtBh7LHDWWrguN
rMSchaiVfibdlSVShoqssnfZOUdw2NeDYzSlZ3+EkiSpsAdHMtJb8LzJs2n//P3SXJaYbmGDt/99
N9KJg0HaV20iYwbSZFabOn8yCg6kmuHq+VtFCzCUxfSiaUEdGofD4LaDuTh3gEG3CmUezg65+DgO
mJXJG4D+y4TBZ+ko6z7d2Z6OohfhsZQh8/UoRUuiJM9Pca/L/Rq22hnO2zJWnYg6LA6Rtxu3bRmo
T3XHy6B+qbTrDcs7BDe+feafN1nO+aVyQaaxak1y0jFtYpqNnJbKTPW4YWIIX/vzVsaHm+if7Vtu
VO5zhnDi1xG/zcbK28dDpB27l5KmgVXF9Q5ECDoo/yTL3DLGXiTV/XmRqyQ/GB+elj03w0jjCIDF
r/uLAwpxybM8e0NfICnurcQBaFlbRpHHtzwqRReYwfkOVfRKMT1pMk9M2LYWJ+A/OoMMpZrbcyOh
IJ6azF1bJVrThZlqS7u0sQdFaOhTJg5RZgyvvQDlOaG9ijPcPt73LQccbw0Gl3gwmAvKL/9fZTNx
e4hMeu5ZeV7fqZO2xJA3lIupudTjSdomqiDD1z0kJAdoleav4CYMe6CzGbcETcos/Q+3CTvTJKDV
xuxTeoszkSIs2wnjLdg9RMn4Eti02FZY//V6cBmZETbA5S/obzD+h89luokmTCkoR5nva/D69S9t
LzF9frDElXO5zXO/0e1G9FPN5sJsLIqNXgYkccjXkGIISiLjsrRyw6W3aS0ywLItS0JLS4HrwDWl
l8lUvLRPbCnDVJfEJuQlqXMITrQmbvNRujKXMNWbDPO3LpGUF/u8j2brjmAby2fifb4G9beg79AQ
jV7sCs2N8np3KczQbKeLFGa8rhjS26KkM00TR51T75bxj92bf7FXmi39TjJ4ULyio77jf6ZBE/q6
lh57XJq1BjQXty46fHdb+8NyzMj1fWw/N59EllcqT2l/5dq83GV+ulDQQY42P93Q+2yCd7fxjyuC
vATGdpzKEjv8V1zmGXMI9LlDrUdwqsdhLlvPm92F8zgfFgDF0ZwaJ54whecmq/8DSh5AnL04YgW5
3i5XmevwVGSgwpuN76h3HMWxSr6WcPFJv9bKgOv35RPXukqup63osgxiOAqQgMDWdbLZTEqkZcMp
2il4hexdeEukytjOhE/tBi1+7MBPFGCFpa/2wo+h2QH7meRKwOLMgG2jd1LcEoTYXCN6OX4setsL
eAIm+mLbLQJ8MZToTbRzI+AWcNJdjdFfj/uSaP3GysU1XrEzShJRBmf2MeGODimw6cEtWhOSgfr8
vPqK5HMKOZeW4zyIjU+SkTEGZW8XcL+P23Yv/C0YAYR2/i1MOS59BP3jvb15MiXQ4WDn7lo1Vqr/
/q5Yhhn/6OY4GHMirFfmRlI0XC9bgLu7C+LlxR4XaJCtpYVdfq8kBBek0MCCIv7/xr7vaRnSDzQD
Cque4N7ClTRhfjmfNQBZVtZQGSxc1vZ7rilfMDt8f6kZ1b/qSrrNFWFj/6nlp2vW9VYlcMKpZ/2+
WEs9c/xSA1tuR7PmsGrfcSTjnUQST0s4588VF0GLOoOIGb4U88tDo6/G0WE4qFYxlmLT6c3UNw8u
9lVChjNh1cvp9VUL/uOZxF0klbTnrHlu0KFsyA2CQ7nxcOH2Ntf35FKM6gMXsFXJ3AJ0yveARPid
IAfYSaNdR55pXp8AsR3VUraKpfwjdQUwLBO87/eYYpTzwRu4oT3fCUhA7KXntQVNc3TwfiwnDpQP
gvWq6ci17ajvH/iM2y7Lp7DXqVBDlpLopVF5FRWMBOJUAHvfLIjL5tt4QCt8e2Le/YIaucFCjjhC
ap7SKutVFmX8Y92gFRc1E+6fqMSbfNRPLa+PevkXQMWKCRQqNFHcDub8D2Tatn9tF+Th0m2usQTk
EUKj0Hd3HrB0SmvZ7Q3LcXkskTfRkTLMVsGcS/N81PrbDT8BIWVHCVg9/JogmAGCn3uayoGN33VM
NxR3XyckeV/9YMPsMc7V+XTDm4jnPKyqjr7VXPabwJN2apiT3+R5LruS5PdwmTotmE6cxm0DMfBU
m0MGHlyOR6FXLpIalPhi7mMu+v34gzWtRKjPaaF91boFU4tJ3F9NNmLiXt7vIH4ga5I8fM99CwIv
1dWlrL4n45cJlEyD6qHWwwzhTPQHntZyARymBK9MQ/m+B/1gy74ebwiFFvUb0ZuKAvhL9GEJJTyw
LMB6B8vkvKTf/XhnZRD108mkCucSZZTcoRjC/4sSSDit1H5O+PSfd0019q6q9nTYZZYyFQmGQmf3
udrvh44ftWFdcT95MQ/gAiF10Ohbn8WbWsCM60fmkLGmZzEnioLliOeDw9T3IWiYfn8cwkQ2GGUt
VSSNdFHVGxOVVIVFsKJWh2+Id3cXJDs/e1caY3RC+V2Zt0jqGIzDSPGn0gIAYcQIrNQCWmwF150+
ySvieCLea2oYJjLKtxu1r5PPumVCq34xBMcpdoPemgolD+dCq6p7RL0MkTC4FIiJ2JH1OBX5gOSx
1+/ORNQUkBsXKW3UepWc3qqvO7o+8xfMu0fYalGMIX3cjMGTCHihOv78tEM/LkVZoG/QWditX/ZK
363mI7Ira/l8/SAoc8xGpULQ5u1lOwNbk6yOWlzJdqfBUxMwG3vKOglgD5s+2YOUYCu8Z74oBv0A
mgyjkmaBPkl7e8m/CYLClPfmhAVGDlwMSNMeGffPxxTyS/NUXSNh9D9Ustdi6gk3gufA8V5oMPnJ
hi8ZUbBE7VQDYiswGzx8rHAnyC7nkAO0gYKC4WN2rChUKGsAqnxFhYzfn13cxhHSPkV+XXaM2DuR
qDPw2oKfl004hq4TEp4owPmYZ79F9B2U4zC2dCLAd3UtGApg2NGVrCOFXbePxSha1gLJAqocavTL
uPakmEJtifMCoXb9VbxyVl+6eUWypwWYvH8VgaCYwdNozpTO08Dh9wPWeQFEf2HFd2BeclJd/pdG
gczT5jfMURyJcKQ6me6NjFSasDYaOTF8I+wANLtEziZHJ//jbRm/unL/JlDgJ5DMZHW4Cy8tNyuE
zFTD4pl+5+T53z59/0T2pDpqBKqjAThsu5V7G6bZ41FwJpa6rb7Hgyx38oVYmG17geuYUJ9IjZu8
KlQlvoccCFd4dI6dsdaeVoTWBmOZqc1gkRmAmYzYi4lMn7chZyFvJfnenS7RJlUqFAlmoyRdmxwr
bCnR4GI2QWw8B9sXWz3H006kFIWNduY6NhckcHxuSXwoBaJa+9HfNwm2tLLtSOQq+/SQQx+E4w1W
zhmugWWkuWBaq/i4jAtsKnfNXd2fMyyWi84xCFIsOQVQz0i0qBd10apyDv+Tjny99b857yR3YrWt
Fg0UJYhAPFGQ2XdgnisT+4ZOYfTRN1JfCNjckcuAXi2f3Bl/SNIvhSVkYysl3c1U3Z3q5D3+ZhAG
vlC8kuxI4mPLM8Sqpyiu22DuJxURSGFmxI/6dC/xMfgouCaYK2wBtsM+e2CNdHA1ueyy7ggeIP9E
RvaMPJdyYvZf1NyFIkCsyF2vkD9kjsJSi4XGU0YdMtvtAWlafx+/aI4xYbO7xkZvKkYeQdplc5c+
qgL8VLYCeEEBRW4I8MZf5B7VJKNlZPUisUZVWjb8QXKAFHqjRoHphHDZdsHpMrASKEpg4t2mRjRl
cMh4G5C10BETYKc6pxkc48KRTNZGgaJShYzmOzSgNTo7IzDjM0PNj5OVSnY47zQG3AApfHCpyoUx
0JiIjNP/B5kCA50m2Xb+nWeadYsdPa6Y7719Bx/4uaE+l0sPEoEnV4IPZUu/WNcINYKcAtHFWXYW
iR68CRCD8L66pmzevqIf3LIl9BVEwi9I5w/cYR6vT128TM9V8kuAXwZjxfozGmrpsVO1P39uXKty
GgzhKhxl7MZyBtaCaZo341/bn8D5XSLNJT89PiGKcsBwYXCTNMx/K+yAxg7kl+YrVSMiIsRqNj+T
zh6Ty8cznLQWEt6blxaNQtcIANmQO5pZeyBtUZXfPDMLWI45CBWfpiyaNJOxhheHyn7EEI68W5YS
+ktimUqhvBriq1O+iRGNxtoiZsXFo6QYj/xjGO5L7iSEqIVMRQ+NJg6Dxo5YxchkGbBR7WYSjw9/
vyQEEMTVrngjMLy/oN3RgY4E10lrk/34yQSSmTitcUjneniWIHlLFFRElKLN+Wx5pxiv9sK8Igky
pw61rmfRJUf/U5nkTfnQqzWRVKRbaCFokQhI6ff67e/bGhKiC/EcndnskUOeR1nQwMdUadyNRCgs
BaFsKLyk2kh03YIfITklCiiupLSPrYDfD2c2f13KwjOFBHGGnQzKhm5sGX54hx0zZN/a+L0fmRKm
B51gqfKL5w9YsYgiYwzsnqdayTio+MR8+mv9Lw5Gf7l/6z1bQ7tVTl2hRMNyzgqPxJpvipMlIafh
Aa6C9qnOXxGOEqGdp2Nakcnx+RoHOKMHmhNbKuz9fRHc1T24GmwALXMFFVq7TI+Tq7CXblD+ine4
0A1M/iFZfBB6+FebMFO7DLXhkmFfnc5C++KajBwsjkQvw/FMgmPKboMVJ2OTgdFTJtP6ZYbXCjhC
lgvcAbvShDyKnN4Y53klSsFtcdIRP2L/0ZE5W3oeu0ZGMyEgxRW5tneoGp+L5BhKkV86R9/m5h8j
78DiPwKYeHSDMIpgmyMU8F7hZcBaguuEYUi+6XNQxyjfCdok2DS1Lm1W159ffy9Oe0yWohQBCGz2
1e5cY9Eq/7LOVFh5Y5rpzRYqP7InROBy9stLLrjSJT7AcMMsOsL9NrKlUWcMn/MSQZcmbyadAyeb
+F50JJn6eo7odCLqSelI82qVgbqtw9m7T/T1BVp9UzSeAVQY7Mk4kbpHy9B4CiEzD/4gMF1ApPq1
5M/zpBd8ZjSz72xGMXAqoZR1/YbkV98GL9UsOjH9hVaMG6o0C1jzw2HTCTqRTHkymC624kjmm/vD
JZVogmC1TlIoVGp+fOeH05OVQFhMqMewaJb1FHGjo4UmVNvpHf8Num81PXXHbH98HomyZek3lYDT
3BoxE2aOT7osHex9t38CcRFg6Uaoo/gwd05tzdU5QB4EKWhy7s2EY0st1Tn+Ua4GWRWDsBO15duQ
bxmTLzdbxtBTVLtnoP5H7mW7wXMiT6GYssLrZ/mPop2gWWVc2YSn8aLoTExzsoRrzFx9fjlvAlF7
kniuADPrClvHKMh7rCKUIhaRuqk6pkqp9tJtfl0MAz8VSsZJANbsMFuN7/j4WxGftiLYRVi4Ed2a
czYuQXwxUkKB8eBolqK4peRF+615suilqPXaJRIfD7duMS+vpgvrZuGtWUfTcHtcBREC+PUwe3ux
eZg26gHMaeKEycLh8uSuGKy9cP1faqP3fLk/emCvbnQQlBT+sKVJSnK24JzapdREAnNYcWFQQFD7
fx5coVSgKjEQFgzV1gVKlGWCIRGlAuzMmKVmy/UpPEXXKeePyCV3ILD6D8CluN7yUjWXDcg5hQrr
L1dkMP7ScMAOnYy0+GADa1pj4POj9fKN2mfgvJL1sT2NIgsRIK9F4038nW3WuDAIm4YtUbDNorwg
AMk3mdFlqGkAmnACNoWJihbS1HqQNbDGgNQBPEwXFQgPMjg7g5c7xlVNiIP2HfJHaQ/KGPeDbSsQ
TllxiGLokg3EV7IVj6IcNbLmydW/I7RzxBdT4QvWurAkcWt58Y1tIA0FJgXCjoXlaVelQ+VxkOhi
zvXJFH8rEDuc2Nj10E1Y/iMRepOFQbr/USEGkjX7ucBQeVaZOwSjUjZxcS9LWLUUgtPNujYIb9L+
PGdt2Y6NwqeOAHzVC/JBQtWUWYIdyz05hzSHdFivb+LF0vXSzgdRViZ8iK6wJV5GP8DRxM8VUNX5
cgvxab6umavDKEG2TQBxsaEkPPEnXyxdIPZjIcptxVCNri5zSJF6qIZ400GV2MOEptn6AWGmel2G
yag9/ZkuRHr1s2Ip35HBKLRL21LVsjNBD/y9Yg+F+sVlX1VA6WpcXqsUzI8qZZjC87njcmcZDPQx
ABgZWydlbjq/c+P11iXbP7kEqqHu2B4AuYDPp/mb6ifIXqysy8r71uTeWPmXsjLOf7ptp9uNqFCk
zIevMb8Asxww6s4I8K0ESReE/ml+1LcVOl0fKTJisaaUlW9PgpwLq3YBpr3b6lQ8TODfMt+XRBGM
+t7EZ4KHQJ6/emODTX+hjJ4ZgPtnoJpQSfTGiaqxsOPEzwI2G0IjG2jc87f5WjWy1KYuucqg4yec
4oIdNxlrW99U1fBK7qkODDdhVS6fo9UQfZRPMA2B69wPfvneVnTJ8wU5kTKfJmfbgaxDEnAcjlyd
1++Z9hjuxUTJK9Mh6G0xUKnXAczs/uQIGa/fz7jbxCHEDI4tkgD+zEhxhvJke2b+JZyVMpEzGHTI
OkAKzzRHaw2cEC0HBdgLsVw1nIVg2a7zhrh5X4Kk4WVXbhgTV2TTbugCsOphtL3o/QvAK5AvAlV1
8w0+d31uqxKZ63NbZHNyGYhu10RXk2bE1mduTs4EBbU4uF/vcnPsrQQfZlnEX43Cjo5jXnHctqqJ
k5JvX58/pyEoK3JzsGRslD+6IE+ASGrf7wpM1vcbA/mqjfcN0sjdwIPreaaypQonJRUmWmw5KHSX
8bR5Dq2PyqyynOA8b0mXQ1PYCMCcTOLXQ6Skm/+QK6WeBv7IE4Ji6yItoWP+W5DxTv1M4Z5cQK5n
Zv6xC4itoU7ZzN++RC8QX2Fx+w+ztxU8Qach2CK56DU97sagRC0ZILz0AeVmIQ/Xoabc4k7gXPHg
TDk9vVA9FN+Hr3JNTjj1w/xmhCVjpDBjW01NyIZ6eE0aXBmoxvE1eqF6WgBjhtxdXDNX1h4NJp/C
9CuXwLkKnAfFUHYhXZSceblXI0KSMZF8yyGtYRc8hPZvFxaOR73Ckv9GlzksESVYgqP0oCOMLAA5
gsn4bHLZCXBtZPeZn7W0wmOiiPB1j43GYQFj4Ac7mA4fxr+KPB6Qw6EreAPgNdC5ZK5GFrno3Bs3
CIKUfGG9m2d7XweP7gyNOuszcOIk3bY/XTDcnMiaaoyFnOB5haD6jg6kaHzKQLY1k0+kQzeH31u5
gbm5y4FJBdWxUu/UO9zhATN9f7H5NlgJw2HcUfIePFFfdLBRlMmVM9+j3QUVVucWbMxwBF/emevT
Z7klXwHRuEKclBqaICOo01u0RDasGyQFeUJ7lzGRJEfCSKg1VR8qLvBmC05IEi7y5fICsiUDT2Tl
hNqQ0mSkn88GpjoD82tVPZ8yB/pVwaxU3oMHpOg2ioBPSCshKJrkw2Xu4Y/3x4zz9Qg7Py1x3o6O
ijw2RpDZgNehySYCEUIFvyVHbgAK2oTG383D48jANn92xpHfggzSFlrEetLJnx/mXnsX/HQc7JOe
xEnzCpjN3zNLcbqn+CdVXe7v21Xbxc9iKaz9uG0WXAXMJNICr0cK8DtjNa/XXOerKslhDPHKeIn0
OXSJ6IusvSP3vT/Cl4DbcuTUPsEE+9QuNhY8KjSx6eGESiwTcmNuc9foIxTHLELymO5BBzzQbGxr
4nfwhZJVzj+rZGTFxiE7VJi8Z49qNVzxaVV7vOda1lKyYCy0gwNvt0dy2LvzRUCUw8m18FddZziS
VOqnRxWy1Mukv6o1TuETFrG3tpqa+AmtJ+ienybLBKaXtVOvqW5OXzwkGzIytek1rwOuUwW4eP7R
Hu7SECwRynJX6bwsC+TnePo4nid0G356AnU/vULmJhNOEPknH24XnMvUIAUM/+925uB0JU6wF3NT
5YtTAXj8GSOHTfRI+QAvXSRWXKvJ2Qy7HBZwtKBenNOUQA5rhm1emaRMrhU3Q9oQ5ghUZcc2x0fb
kb8JZU/P4SmiD1uIDwU6AHLWgVIAnD9UMPEoRjDweBv8k03BdeeC1NS4eiDsSwy6bxmbBNxuyRIY
/Gd04MPQ110jz9Odhm0EJqmiLmUnuNdd3B+r1+sxYJjCyGgT1z+YBvE87GE77PbNSIJx1HOK1HeT
/AwrEgmAowL3jFMnwmsVIvZ5UD/O/U7oFNINv+gFTnokhtpzj/dRqzm224kPXWHHPt7whlZG2jFD
93mJ/Si58q4Ptwskxhrxld/gNbvi81Ba83jIAVloHzUZlw9UX2VI0knAN8z34EeoQOoFexdYOXKO
vMV8sOT8vxFFuCNV4XqaMoWgPxoUD0GDpQU3KoenOqdGK3h0b3mAV3uwRjBBCcUZgtX0bIrRzFGe
0RDfbPKaVe6QdeG4aKsfebs57NrvkVL2Kj4L/5GtWrxMGr9V5z33kLHm8BWD7O02OU9RC6/GUjCk
ncu/UNceUeNwPbfeB0LXWJ0UFtZl9yanR/1dt682VcieHvVDiZe5vfLO+jjV/IHGk6KmHJE7LnjV
kQ7J/2bBDaT2N2b/iqiC2/MXxrmC5Hqg74/r8S3HiLxVS2T+mQPTGfp/KAFHzvdk7PcjXaMKrKOj
tCYB4cpLWRIMwntly3VM2tUH/vTUFCfH6/DkL1CTZVbW1oJU5bbu5ITVg/DkwlorhZYzcoTH81av
las8bam6bAU70inDCewZ2yEQaQEX/EOBTlX3yGZ7uEYQhTfqa1WAxbN03+m9ih2Az/kLIthpLx7o
iJeHXVOAWKGwfC1oBWdGutb8NIIXxriZWPVzT+AYXKMHcb+VidlwjLndyA4wyGRrRAu9QXXD+v3+
QPcptUb7L/7fjm7qEc99l8Ow0auhAeNzkxK/X3dGb4hdxM45zWNdv518gxLMxuTWQ2J6QL/gROTh
KVy1jHu30vjPgxZqm5Ve4M5Tm6hDmTAEUc6bry2fUypMRlYuCJJvcmGwAvcpB8YN8SbnXFTltFGk
sjFiBpyig710gNr7bK3BS7SxNM5iAPY1Dej1whdcl01MI8uLoPKHOtwA+9aFeyGJrfJ+sJnhXFrX
u5e/uR5Iqcdx08GMozN0RtY/CN5To/ucfzCbA8amIs3DJyKbUaBtW+VVaNZOmlrMvUkuTnFMGvB6
8dgKSAsU3cYpc5hm0BH5z8LBqjAsOTVxwbmfVqaZYe6ISQmgSFuZBOXQnK6XR0XX4ff2Saiqi++Z
DYQLWiHrhkQKJfjv3YLjvjWFBEOAcRLNRLuysbevgzBaDPQYfDY+B/cV0qrYHHTPkmwajT7cKxR3
A8P7VH1HssupS1oekYIMpzTM6T524jC4Q6kQ7TN0wEyPavyqyH6FkY0bifoTQUD+Yl5IWt0Ab8aj
viL0NUlryUAlOVUX1ZrofIEt6KJIP5K2kMfqA0YYuYoX3BtnICrT4O2K4lX0s1oh0WtqJCdUZ/Zh
dRfJ1eECL0fKwY+BLgVXW11d/kqBr5cferZCVdIdERu7TbuiTAGLZ8FO9Q+PKyL/de/BJJ0k2aWH
ud3VblJSXdOaCvaEzNQWkyBT87rcUKCwYlZKNAN3D0VCHbANR3Jp98ayJ8bH9DlL+mswo9hl40OS
NLGyeqLPVWUNgdk/6oxJvm87namqyAPQAtLYVRH+y0NpBylqkHOABELmJAy8P8zMhDDuLyHJR2Q+
3Uj0ouOKPIboqZhszHPowXdiYqAXtGGDGF/lOMFK4jRWL8virLCUnmr+HXqVfKMU810BkMYq4oyu
lVdfIFIkA4voCrq+Ms4UwltfHM/9SJ3WJWUMdTfczA8gS21gFUwszVVoStbUtnpn8QeJDgjEvIur
JaymePb7xBNSWXXtbe3SiH1+yRki4otwA7aVhB4NRqM8/wnBUAP1rIHO60igHcuhyf4dA9BVwrCB
+w3Z7ymiKFt7RsXIC/PiuQCKRGZ2wapJuBPGCj75/Np1YoAviOcSiEPBMlniMwqitMq1oB0zQ3DY
KFw7mo0qChyYuKsFlAOi+4pdI2qeaP4wXP2nigOQ/DMUGbxIFNti3evUhbFqEWdEuGs6Ao6CQAO1
ieD0KQTeFhL2S5TwW+PIknCDNz5LHyhCqiQu1+uIH99K/xHKlLixU4IXQIQslu7ucWXc7UV2FOTG
8xXUwGItyh7zGSj7lJbAhsLFv067OGS1W4figuOtLer9y2KOHGkNzj0wix3GkCnj+bOoDsyb3LfH
dYA7CiXWW+HDE9MnW4i+qHUOol8MlNE2T46OWqvH5ZCXhJKEIPL7YnP8tNoI9W8Y4sgMYTDgV1wQ
9g0xVbPuZcy+6MDSWRud8cNMxvfCYnl++WSsJGVMDnxNPVtxQAj6ANVnFXCrllbSMgrpov9YToxC
2a8QXOlCxFU3ulj+OlKek5ZD8Pfhfktdz0I4C58ObIBjIq0xP9aXeqHSfDJvyN5akorIoFS4ijIk
i/SZjHS4r4+nSFLrt4S0hmxw/P17bsGA0vJzyjcoNFsOiXEjP4/5Rmad8aXPvWtQfq38naLOLPsk
31F8DnslMHLcbe4cJkfrEHJB98H57G9Och0LXgZrC/jccsmCgF6rS34Xk/HmBI7gnygQjwMmfwxL
W+EhOl/q3S0pNB32KcFM12FvvQo9xHGN0SOK+5I5VfZWM97S5n9ZK1g867DFdImhHbAIDfsOxuPD
ip2D+N3J8KaB0Z6sUDSqCOUymU5ssKnajrIB12QBzaqSALdd4EVNYkBAEYZoe6Jh1ftJoMgF92/c
mT+GmNUlCeu0fzg0N9xUzEmfRl2Xh8LFC8nXlzjyab4kjnCq6Ypx/kVx4A2fwwbzDCclHJU6tFxn
OeUYx6nkH49mca5lCugzyO65dfGghAKhh63nkIilPHRywcjaMVFZFxYFQbpqKqlaFnjgaXrcIJUh
ePPRHLE1xBsuzlCppl5ILVEQ+nHSG3E52wycukCjDD41YlejK2+r02/AwSH/sRUPVrnwds7V+zSv
nbL6HuRaq8z4Eih+5VV9SjLUqt/QqE5acY3QMItilYXTjEiM4GC0VJaCukFaLrcQ56RA/M6RxIlN
9Y9oKq42lZfU38LBhWKY1bbDBq5lvncnQ4S9rdlD6u5tfdFZ6TTDmsVFjv5lLIVLWgFbJ/MT/xOW
dAiNa/2rXIfQeGgO8fZ0Hu5SX6pkf6pnRqCmq0FNI1X0SSmV5w5s7lucHZoxSB78S3DbfMahghAS
w9qOkm7FlSedg7+G40EtE/v17dWEVGZm56j8b9fvz9Ublc3XrXdn17xnqa7vi+hveX4yRoth0Li8
nOq7IT3bW8f7AdkWplu6poq5GKaG6eA1eXzZqsupCEDEddVBhsVwF8/VGNIzIKqipgpJ1EAytkYf
1IOwm2052AjcAAYrURyfnkeoFM0smB1bzUmmJuHPCY4MpclZqG4D5x1xnqaMeHgnCydgt59oL4M8
E4lx7zqSyRkAqxAAxghVTx30X53BKN8ugGn9HX0pRDoOOG9fxSBeurm71qowFyYhDgo2j0FP/Pla
EEhFABiEynzp8dYTSpaoPEWeHkGGGUqaSvVxp8IPHP9I4h80pyqpcD2RDM2/dsq+sUiK5yXNDL46
eeZDdPvufkP/qp3m61rbsidVfUB2zo4rXkZb746YG/mF8U1oXyO0SPESVoXNIqgRqI7wl6EOVGj7
rW0p7ComYSP5xO2gZr+rrpnEV3sDEgwbUrFqMppvJh77CZl3ghKni9AjUXcGo6yFIBP+GDpK7obr
tuYiB7j3UXdiPzxEdWJeqKB9/X5fXQ3pJcmXSRoZyEAUsfiaUssulGPz5iK0vd4G3Icyr9T/8Uba
vaNLXmwsYsGlGrGZyOiAcoaHABAs/DGwvMpAF710d+xFiTVZz/NqQqrkDv1/7IfcIk649jzwxp+U
If2kZkVW+mELRucyabmyAo4wDZnVDP2FoEc7NeY/hDFDsCpJpVrbbumTJr8Q0qn0GNgW2SRsWwEE
Ta6WOJbaSHysoTIkD0kNc5LO64rSaIE3hgdPXZoPdisNpSWXPRSksXx3m+kyxQLk9HYfWHsg/p/L
i/iqLqWGklzPFGp+pPjy/TOASbgvNEdkF5tLkrXwREpf7ytch1SKczCzbcJg9UhtZdxBE80eSxKK
D3jEtoHzDKHxedtDaZphrDUGWJwPW88r7b+44VbnKUVfhjRBroe1ss7S0rxpS29721IwxdxMBWJh
4zMQcMOf1iSTKsAqlnymIa29m8s/ST/3YJEyvzVRqrvRnaVLVNAo9m1/OXuoQXzl5Rp0ZkgYWu3H
5wkCucppyTAxX4bsq7BeW5dMuqqR46on8lzfZcGxEDNteRKHvcYinpmqUUaCmdCalQ1BQOs1rzbh
G8SIM20lCkmckNfVVnWnPcQXH9HN7Lv+vE0CQUoASpCcjz2VF3YCVpIClIGGl6jmk7lRmNpoEzRZ
qEqbAcGuDvJZKVf7oDmustXMAmehfSTNKPVCuEf4eh/67dP7Nx8mU9jv13JvXSPDss39nQXThh8U
r7gviegFmm5qbnDUpj68H8H6CaoK80KK9ucNbvdKQcnexvUC/GEbZz/Ja2H+MVNV/3ufGRqWiU/6
DrubiIZ1Ft/+Q8hQkQOrJZZ4ZCIM17zohp0CvUJEf2O+6IRKL78Mf2yJ3tu9SFmdyp/eYZsV7QD6
lMtTOTto8hwZRa2YTdtR5GmDS0SWBGJyklNXUcRGaGA5rXe+shFimELV41Pd0TCQvcHaLvFTmuYY
UdcK89ik/cnXuMejDuQW5hHcE9+MnBFx8wIR15Udv42Hk6UTdkZrYmK+e++zXwAAo77nhNuU6WQ/
WZbWceKsOKaLkiwPw2R6C2SAbf2aYOnYi0lqCQ6yPqJ0p8RImiWH1DgGW068GhxZn4Pu9idWXDb6
a0ADFLsS4UIa9hZcjzG45+RNBEgK04/jbfR+TVWfG89cJG7kLva4rKgxGqmMrD69+iL8Ok7ygHN9
d3muwI/gjPb5O3qsi/Rj7xaGW34EzjVA6AK/C8Ru9ZFMbTNmAkIwRD/H986UfdgvFfcFlAtRw6lX
NpsiFiqnXllvevClGAqyqxMKw6ZQeAonN6PMbzujY3ex87hpQOu1Cd62DjRox9tOVFY0WEXJWzPH
wco3ACv/q+ICcSM4WclE3m52oEKEGBO9C4iglyzqo7rQRVGnurUzpKE43pqdk3v2fK2ApYUTmIiy
oRCWkYuOsh5HeDHvxt875uxiqVIPcs+VRxUOrnrbn8beyI6oKsTxnEjnJsh5O7ei71VCjOTF15lu
4Qc4h/wEYuhFJR5isQyXsKCco4tTKZIF0X9KhZ4qhMnKgPrUSFK3aqdiI9T6X65kMudWFKwXhRcr
6vKIhcHhAFpQosBEJ5VLQDDFMcJjI8edhkXw2/5GEsYU8J4Gqep3xV6kvWQj38nLjF6px6hXO6FV
BIbfsM5woSX/fHBMt+/PLoZEFjmQ/eMBcDTRe9ZOR92ybM8dRNL5N0fm+jlKKxoUEDpX/ut2hMBU
9NV1zGdWfKUK15j5LUK5OopZiscDPXOIQlq9uJBJegR4CfVYxvijYuyKhq33E/ZbbrpWVArowDxS
lj7yJaP5HetPt/sO66h4N5smjztzen8wiWMA2tUPunUusAyL7UowiYeNHgp5aa0VChGIw55LCtj5
94c7qBStfr6kytwfDLREodLpDOwx0sAz/eFaMTsD3HR67+Kek7rKj5vRttMZbBgF7XZbagt7A/rX
XlGW9qx+ulHkd5kLE2o+e3JvYHnvXhHs0/xeGEwVl2ONr8n7LYgRXVT7WmbfB9+vUaZJOVFebvBa
dyDnhjBk57Pw3NfxKWiFtp5tbCmVVS7N350bsz1r+r44JEGEL7tuF0L092OE9+p3rcfTkgNG8lXr
ISyYWYFPRxNqPNJr880pHDM8JknhwzdEQ7bmBAtgt/jTj4x3NmX554e3cK0Ir+Ps/uJHbRiSGu1e
Gp6ZlNjP0scsJIuXGPOTvXEXEpdn4bQ/8NQbMvILkhQvz8Y3Td/84W4f/RGipPBzZphs7TNgaHzM
4qfwcNwirLbl3wJY/tk85pTDnmcWAx1afuec+Nj6mxWybU+06fJNo/rIluyJ6x1QbyspgAce8Fyq
pkOZF2thyhE4Qgpjui8ui0ISNcOq6OKJkQNG18A5DarvWS67UXCtrFB58+ynn+AeFQCFxlehG6Fg
zFnVbfyYB81FwCrTPw3dWhiCtxxUkMqbYnzHtc/3l4nBDR+KRlJhl+M572TzWo0MkDr5Z5CO99dp
XOJHrHx6FnMBCe9CAPbYh9DVTfqO0cpxlj2Yldcad4fGQYfYycLjG8eLkllAEc7+VwdBUecUL3WM
QYZY8ZzQB59VlhhEWSmQGDxX3vodvRpU7CjCsxXtu9NDvYVSNmu5Ew9cnmThIIPYoOJeeXj6nQIU
ZGvZ0vaA0RQB16nEYrFEnK9G3H+vZnPB1RmI+MiHz9yeNT5LX3uK/cFaVEPPJKzVGfRiJOKiyCtZ
kgT9RAWget+BHKt4ipJd/Ww7WubAbQ7b68pj8WiaT8HaKKXaY/R3MpfN/vWOC307K8SBRZXMhauO
DslSmwKmev3s0xtEl3sWavBaWYzp6P1+VkiH5uE8TWuUImQVvSO0V4H0DFIXmTgmUi3p+ezI0IGX
0rJdBR53Wh79DsH7qnEJdfhzdLiaecFXnRLpOR1e4nhtt+EuAAa+YbwL0gHiFWmHLx9aEjTKGJOV
VXZRtaI2rJd8lvARjRXorCXhZ3znbJoZMb8jCRKEztTH9Pvp7wu5467uUIEA33q4z02c2HlUhSE9
ANdlKzCoGrrhXiSYJyY2a+0WcV/+SlEnYliGml6FvaiWaJ4CoQ+Y5fXx6hfl/DoCGmMqvMdeOraK
FO80kwwcQDgTKiHmGdNxVJAUHFT7S9jkdiDKk/BFhBwJrjmnc31Df2jYsCzLNVZlL/LuJG4152C4
Ers29PeDEi4qUvXpQTEvbsQQ8fsGaFYL6m50fF3MSBPb5ZTMHzm5rxoB7DhNr9DxE+rQTL4YWs5q
9+49CCO3tAXj9Ok1wKqP5mlDqUPy+chCp9LqTlkNfaB3V1yEbr6QmtRTdcBtsUpK5l56iNOAHZZ1
5MaQemMlhOK56A6ARIgEnIeyb04LFfkA606zEXv0mjAd6EReZid25+d9nLEfGaMuS/jxzz5yTPTo
TiLccm7TURmqr5ygBPuGsEFjavoPx6GGlHaOWrsmNfSpuQKxEKJPdLEz7jQJN/0zXBm6FtpNmygH
UmjC0KRdwgTsXKx2BKeOCBX39Q46X1KGYKUzcbsSUfGNxT12DGTVexXllxeHtJDGllLKnGOIbfre
bFhfplvhavwXbVVlXceiG/4KDTJVIFRJmSVEEO/44+H9PSf1ne+AoK9pC72pH9k/OwlBLVwPRSq9
flPTeCyG1YRI7S7mHWBe5AXQznkJEU+cLOHq8X+dIgYct5Wi9CC9S2coa256XS1fOJh2Yy9q/sgv
TWNzOEAWrdfBKpmPN1Hthrbeerj2bpXABP0eltUBUtTHEyr65juvgoKsqKg0JCmr4H7OjMfpIB2L
Yivsx2wd2oo53/4TbPb1ZnWNbB7GvpFlDIOCkRjKbUyjLcTMmv00xk015gkMi0SfNbQDzwLfngrX
q7IySSkGFDJQde/qF7csl5aM1J4QIijkcV4Rh0V9W712I2Hl+XDbftdkuC5BpqfPObRb5QzDgcPX
trOzURtizDkqefJQTgEuZnvHApDzN6dN2756gA+1hadApTEB1SPL4kLxyeN2MUtAaX+40LPBXPlG
g9l7PNBaTNSxU7yV9wGD9tV5JUJrZNABxZwG9fsI7hgNLAyr4MP1pNeW7b3QIcBQlvQ5H4kXStp7
oWU2/MHAqHaasIhI/y1QqqYYQeczzeurIldSPBb4CFI73izRueKYIwOwW+BMKGyp+cbzBwFkvRCH
e9Q8KNIibYX4gXLt0pax87WzaaWvkK/6ztPhTIyPPyJd496dX3J3erEIjkq71ReOij3QdT4cTAPj
x6QaRVVl/hwen24pW0gPOIDePP3BhZVir9adz4ATjb/k4XilePMJ5yL5d777Quv783StiIn5n/mu
oEZMFF+SkH50ritgh00fhbSI8kgRQi6Ik6vWKFLNJqGCh1U3VVHh16M1Cbz2IOOlKJ2YnWtwyuNX
zKwS8zmR4gw2fxxdJANSFAzQ7QL/VFa69GS7SNObvGjSk7fQ9ZGFm+Xcwsc5DZxni4LrQ26NhPi7
P9N+yotsb1xJcIvF6tZsvz6g4sIg44ZRTMGmebhMnFhOiSIDeMmDKqqfU8g+qNhi506pbjhn3NKQ
QQDjh+5ZfWqj1iJLokKlzoWwDTa/xD4txlgWlgKgVP79ksq9uZyfPMzSpr32AfC+YYGrJV1sXr4N
hk2Zg1cVMLpZlvDLlzj7RDzZHwitJrHUHtd4XHU9NibaC2QxK8gdMME4Fz1pVuCg8Sp2ooep0EYh
VHC68TqqDHaydmJjtGIYhY08A908+EecT6k4B+cwmKXcVKaTo6YehMWwgWLTbEtxDnr9HyZf68cq
dLJN9isxpys42Xy5zHRFl6daf2SqoLGUCq6GzOh4paI6m71skCdj24sg7yU2Shvc32C+PTGo3NI9
ksTkZeZfO5OldXWYAAtBxWbSIFWn0sPNItCvKCAEOB1ez2CfUh+fE3BVv6JYokNE6rYmPPNzWsov
VJ66BFD7O5Ub3X9ukoCF5xJa60MdcHhPsRC18pHCMvv251c79VcC/OxFrnrD7tn173ydK3IREE2d
OAUQsUWEuSKaYi6U66J70K0J/7yaE9o/5x7kYYIAvOOnN7T36hJ6Km0+6OgkTJZEcfW8dQmQR4/p
Ve7XyATWX9X2SCgJpVYTrc7UWbvltTzv+SYFfjOM8AitfkzBW30TuLZe7f6Mjz8qZN315SiML+qG
OL6jF5Gj33NStTxcAz5H9zVP3ALm6METwJxcLI9/PCh5AbibhPuZFWrjLGbvJLlqdITNv989TI8Z
qjpcgxbtG8sJnoP24DfB3Xeqa8NKJNm37qYof6wgCtoBtHQNWbh2hr9Xuzz/yKpY69RpJy4f58RG
zAw1BTM/GDDT3W8SI3ifF2arU4QCCXflbiwomXxah106GQZ0q1NnD93lVNKKI7wxaxHnMA7Rvh2J
IXHMhboVS3eEomYH6/1PcaCsA4kfBNTb2wnZauGhxphHixiAIyqDYJwWY6wxHY+Y2v6wlc6tzeCr
Ud4Ypv1MZvB5DCgr0lcHpjIuw+gOgMSP7NH9apdlWNLuN274pXJi87Tfk2LHiSLFc8l6QO9SuKtS
F5kpgDvq6fnkObmqz2FAx5FE0bMWpHHZ25FLtkjhaFNoyE3rP4MOW+wl99CxxPYlx0xyYjL3CQNr
6RyCM/3KaNnPGFqXVgAaa4lVddrc0RZV/oDkf6nq0AE/bPCJXtFgFchTnDR3D+2f1+N3JQuA8Bj9
w5PBoCZVF2xYvKltmRT2FSkgHZ6Mi0CgS9QLIT5OBIFJ/38wbJ4v84Fo8YeYemJyaYplPRCIm5mE
NhYXHhGgnIA/rZlEiPYxDhWdlW7MSqxkGlFhrDbe6s2zRiwCHzhqrgEt3IShvY+/nY3WALaYCHZt
r98b+1Z5TG4YNGQzF/k7bsNcQGA3Afh0166ZAeAuVq1UroRVdz6aeUEpj02Zc6IVH/LiDBeeU61g
pfMd3OhLOCAzHJDT4vxOWq+3xa0zR2Xl+CoRwZgO+RyNF18b3l/enPv7NOcXMzmI/Fi/4ionfwLp
mMDRDEhW1Rrhmm40DN7oxUp2Bhhk0QtLvVLlsfxMDYzHt/C3GMHrL+CqcwAPX3aRyYcNILlJmuDe
IQeNY6Zc3MqPXBgDVt+Tz14m/jEuRb3usqYRgmHdpqXlAaCbOmuJGZxaiVhme9IHcBQ88R6NDEvQ
rkhpIukLx3M6toOlrV8I0IOQZWiZ7tflZbGWaVqx8zmrGfg9efGKA/DgZ79kMk6Oo93+TqBo8tEk
Ps6pcj+uL31sV43mPL16s7liaBTH+qhXMZgHoBPpuL3an5khIWa7zE/+4ACoDRO6NmbKyh92xv3b
U7BomeyWmJfjr0cZspuhMRvpMnyW6/I+KlDuk6/Aowawg9f/s0N+DvHFRlkSQhZ59JuxfreDJY62
TcSU8bWiuUhsSfhODW5U5QL/RpBGk1jCcr5rlaGOjWY4noa1QrV31LN5m/NKFQvoZilnhHl8qRmR
RNndmURPMsmIwmWgb+t1a/mKox8kO+aLipxi/e4axqMtmt6IO8Eais/axqmKf25xWD0vfHLStK1d
jIES+KZzNb0/1051TOXSRB0LvrKJWg8PiwYnjqo+UVhk6SRR/9et/9dFMR1os3dILYEKQhLSt0lm
/6DGi2h2WdNr+mdMVk6KEGeHiUtrvAV+MR1yvt56YEpa5BuX0D2fkvSPPLb4cUoKCgBIQSSCfIAh
qnPuslQI9wFpAOv9h4jXdHzN+Zf0mDTERh+z0rZJExpoPTq7SVphQnIVCbHkfWUMH24jPXwWWnir
avdDManCoU0CMdvDBcAGKgUatuENqW/ZlTMLkgLC9ido+U3UKtKWae86ocw+o7o23DYFz5TmXTHY
0C2hFNKJVgYfTvI8lbxnMqIFEUUtFELyWNFIwL7fbGHKUWHXde1Jqlx50u/C/FydfE2Oosg0IVf/
iRezA9bekDYCynqz1zmuhySdh9Lxya8vnfnQss8bPZPIxT95xJNSCPALSC9X10K0tCIfRSWUGsFJ
2/aGvRjLnVbZHhhDgsluS2D5aCxGYU8ERb4bK0jXpXfNOoo62LfsedxZr/6ICnUKCXkbPjL7xM63
7MkbjUfbzoOgYGZPdUGU8iwVYUK+QJukaK5haQ0kZ1MTIAPWnAQk+Qsyhjz5CVGkyZjeFvPdUrIK
/bciNbOqwEixwiO/tV4W/aeCkHFIjn9CGJtX/L1evWUKK2XteHEkZVpHZae5jVH8nM9LTuQqH2a4
3tJg545Baq8+KMDSYOS/MawARK9uW241I9mVlReBGtrmJMTLTsvnplMqtmFqcNFULLOgWhp1lcSI
i58MNqicJ2hcBMvl1A+pHvA0YAfZI0TcZDIHkAOvtSPWbCiqzKNjjT3JKw9z1E7Cq+CEYZfIzt8Z
6cZKquf++e19FRMjPDNKhLZYjre86UmVO6HAhrJHSZcetieCRsEjF/4psa2Z0gRzEXh7yi+ECIQg
fK1WKeuqG1hszoK7zo7fmceJXyl1ugPe3SAMJF9Mvwcik8B2n/TKG3hGveI7B/k3HtVps24osbcU
V0W8X1CQF3DIXwi4RhopWji0WhL/vNFhOd3eFWoRzI/GhVQIdqOYGxs9ukplAaFioH0jzTbYVjJ5
F2DYdU7sXnRMPJA23IA+XlTHafB3sSxkw9AbTewct+LVqIle9vX9nJsXTLvlzRdrx6fM9Qtxbxck
31Gx6SjJUeifmrTIqE0VEe54HjOozxGwOTkraEkI46RNA6U+IIl9UNXE+ocG34ZEW+BrCHwP6Dq0
xP9azDemkrOw0kHv/dpYqWBFn8l5ZrYL6hWeZbNkehabCZEdz81flrS+WTU2L0DCqiJ6OUAaHRNJ
CcgH80Ja+V8Dpglu4SUKB0AFKbcoiJj5p7hvsnYZ/zcVXvG+LBY2XUqaPTTHBHKliGD1xjfKMhTS
LxyALKH0xAuqoY8LjGjSZcNxDlFqYqWZ7ofU2xaMjMeCQ7yT6uGs61ghcO1Ym77GM52NE2/+TIcp
L9m0c9ER5Le3T+uhSj97k8m7lfqws9/rqP5J9ESQ3bjprh/lREFn+6rUevh8KFfczmXomZVxmc3Q
886aUFAX1Rk6Ywz0xDspfpdld/5BGYnSb+mCPg3cCO1iV/w2+Fl2vsYwdFkqNki34C+o8z64H/FS
Z5JpYkIsasV1pmSHBVmkhcSQE0Iv2vgeoPmG+xL+40zbfQeePc2Txr9HTHMBJXwlxSRG8F8l5ku6
yH9oWo1aTQ1AuN9k107AzerNxl/1+OjTXMvQTTojq6BxbyaeL/JxZnwbvnCr+u1jAuT77gYvjN/s
QsfFrO2jfg5pwuVak/eqi3tKF7pw1KQExZ5fjrBLwzO+cUHWVTnCzmTBe5XQt3OLAmxDqqf3j1+c
2YBdj67K/IbB0UyryP8aX9Bylxp49JtfibpyGDZPLolspZDba8WcYwQqXxuVhR/hEJDnMdbgc8rM
a6YznWIv1N3vg97KoH0Du8INg2fVwIA0LIkk3MyY4ae1fSPQD7fqXWbX54ifOT+8ebKtKSQhq5I6
O/oFHJXhRsBrY9yoqeih8Hj/80GsWvqwEZRGi7z/QX5nUYF0ThKQGgR1qWYmvUybhP1lQ7hN5Vw0
+G0ve4SxIBzWgekXIEU4S0ox9gs4kYm2IgVVtUxeC6QU73ggWnIFQ6CzlhHBc9KHThtvPfPMvJG8
dJyadlPvk6WNZTExTXoIWVxNnys4tzl1BxIgxNk9IRmd0hdIpVeEtQSecfg7klzJpA9y70eprbUK
t6X5Fm3FPMwMLNYWLsyytugthETrNlgaMJik94oeHONqP21/7Sc39HSjd2QhpA6VGAbClJeFIIfz
2i/OeiTzKnsiZsRcDt1fFcHnvYopSy2QGoZF2yJnk2tzBpqLpyKPGAseQu3MMdOSJTlrQorNeF4+
DP5/lvT25nB+Iq3Rd6X7abimh13YtizVlc58UGTrfzox0EwS4nZKCdm2l+lMN0k0G7FaKds54T4d
2kEMIzFwf9cSBmZfWNx48tITSBtzGC69kZ3fGljcXB2qfjhIIUwBuwM8UvevbIlNiIzNZdMKXOO5
P7I9Om+NQMIO2y59kpkWvs0tIDazsQD0ushR8pox8aU5v227Fxjg0RW4kHugKB4AZFxKFa1cdpAO
nlY6f3y2LyrVugz223KQ4MaidlSL/rM+4u9J48TQuz4xpCLcMh0Rwt7OlMbeuQJZvmCcyyK7kbGr
+unTaQSjr4wVq/zQ1GZCrU1tm/5RMeo2O86e666hcnfDotlzkR3uulOc/B93sD9XrI9YolGYlMVr
gM0va1dFJuLZg5rct2S4dWSwp62OL2MdiyZJgBkHbGBXzYBqUF8JfwqbbfqOFJdEZKIxSs4JOrwb
5kjsIcMMdqANIARqR+DBER29uDMOrCPhf3VAabdzyydePpaUdf6svBoIidqotNoMkXB+wQ10zwba
NDdZ4wO9+F52/s2xr9FB1YqwtasALi/IaHb6UKdTeuUOjuJvu8B6nzDNHuHkz949q/u/K87VbehD
kxfVda+H0N3hbhbNJVtFZR/UQAQ1UZRgvQpWl9A3gSXZQF8q0g5kX1si3FtAxs71GfieRJFCalq5
cIBWyJ4Q4EeMVPyKd4zklQOMs+6ex+y6qo8MrA+iqkI2mv+Ltu/IfYlO05L+BUkEvV40y5DaGXCc
dPbH7vQzOYkayELyK2TF/tM3jZUQAOwt0ADgCNnBO8Ubx9NJhZALLQTZBQ4fCPPn3GyJCM7fS/y/
iTtQMUr6FKmKwW6iRj+6DsELmx7pwgoly20bXjMvRRs+j7nAZkgybe2sdMyHe2jnP3LUXmjGVGvd
nnWTVLrbjjNdkSxGkHwzW3YgVfN6hDdGnvsvuW2koMvdC3u6gu0YUEOPX69+pMGDK6gf9QqBFMLI
9I2nR4EcWTKSlx8nf/akO9rHDGw1Ie4ZIinMinvdHDoVN+dFQLXxBF3B/ss75OYwaF2MUSO2BBIX
j7qYoIMyfY5RakuEFIOeKP5Ir/3ib2cb5IlaWFMDfBOWUWMYwrY1Tr3hEn3yf0FL+2ooTdfTFBBy
OQX/6ozCfNDumy+8T1yygR48nVz7zH6U01pgs7xF13GQxx9hbmt/asOqS0EYzRSJkLaVvy+94XJZ
GFKmntoiLNyNRNMs85nm/eWeTq9ppEFYv/+YjpDQyY8PXat61+9A5ObBfL/UWSrXnjlg2ncY9LOh
PVRtlD05WN+ZDAgpzb8LGHGcDWgeMjFLjOVfY9Jl8MgiPaWg/tf246dtWdyS/BcFj/UGS3j5UNTL
bx/cRWH2XScHCZfFeuvzJQI4MJ6sm6pa9KXlHr0Job8792yoeEulq2ur98qbArlEqMDKtzk2yw8+
JTL0E6+iTmB7dmQtgxZ5Jr2MFeg9uyrWSO6qWHrHcDNrI8Bs+taTJhAnPE8IrIJkbEoSnWVWUw5I
VyFA0SwcF46BcxYcNoqFxStk3XRpW9WrnTzvYYJ7AQ4hABpX04GU7brQnS06D2VSfGsh+IurpWw/
hBpF0AFwe6uKtDm7euPqW+ZqvNcwfneqQgKBQKDS7zoLhIll7AF7/xiElYJLasdzPpbqkcXSMeX1
3SoptWhC21yCow5va0D5fao97qFFfwt08zT8YnEHrm5B7u9reeVLC7XvQC83t0Hh4UdXLvxear1+
WKrbyoI4EUUJIdibrLkHjUb1LkB+1aUE7Y1sPTdK6LPraMEIbwrutjEDubEXCGHS89PNHLJlpU1X
HOFpHN2BVSQSquJoMMYNV72It36RmwCu3eFPH46jYPzzD7tPP0W8z41pAyIRPVKnjfvPj5fkbeSC
DJL+cRX1gD8a2woCYVVl56htD3sQkNSoa86CUisjvKYUVbTuX5/m/d86IiU+5wxDAv/C94KiuhdO
QKuvFqyuafQPPkNBxoFIn6LR36MNKLFPJ4tXDePB5UV+iA6w7le5hQ6pWWCVnDEye+Ox06b1VGt7
h6CC6BMXM8moQuuH4cH1WyCjEd7tHZ2QJYn+bMqh2lC4a52yjlILvJuWt3vR1uL6DqOvo5bmjmom
OxcUnextPKE560ZdBCyHYWWSu1bJUSDYItbqHJR/MnWFyu9y7tGlIa0Rlr3dj3+ffKfDvSmq87wH
GfURCvdpfc3q17u1F57PLzJrgoy2Q9h2OUmfkLl1s7bzm0NbgeCP7DE2m1XpMBNnsSomjbbXzEqS
Y7bQ//DxvC3RGTRZoiaSt4r88ohVWGoUcFba8fe0LQ+km9KLWqDpoP7ag3062+6NxIKy7wExvESI
bLuS921KESbV2wsoKf8TylPA3zRSme0GSmB6ckSp7SAGrRc9P6ImiQ9hq3HqlMhjBe2qwhoJjuS0
JDFF/lYGHDCbyZpdesFLdb0/QLPtVHIrYYt6VmpN0C/Uyi2/rE6U9aJiEFxOsNlZEAyUm4phKBkb
R6LGuUaCjQ9K1eCntilqY0VvZluvaIGMjGRSDjptMRljc1xkvLSrUylySY9Gv1yR7pKFi2FBcF9s
P1/itff5pqZjrQiwj0KZdHkM2mrAD3JokrNJWfmQdnKLtLJtkU20ALqBfHZMCDOitlQS17A6uXrA
8bQZYMkx5OwjwkNTKBwxOaWgmjrd5ETQOaL5q2i9MGir3SRwxsbRfBanJQYoi9ktE+CU9PUOMjNm
VtPMxKM4NenCVd5OU20vGPwV5hgUi9FExGQWJ6BBBld4TVJoqjzVicK5hMrsspHc4ZMPCOE5BKrc
t6TgfayZbH6/RgymGw1tGFipXYQ9MrlPm8H3nPEwjB0UhEOK1Aq4rFW0lbehDXLyxHPExVRW0UBo
Y6zKHOmowMDY6gC3N0DERf2+rzuQnrV8gGhVoT99gt1Sa4AuvInhK7NvBaZo+HbYI2FIyinL980s
FIKUykmlujteNqEN821ILTi+FXm7lxTOrxl63JmwCqdSLK3fI5VES1Ev5Ux2Quz6MCFelaYp8LJo
wrjlaaJnBG6GobkMNzU42TnUPilHfrJn5vLTs5OTwmIGvAlEfdiy8H6m58PMO2Io6Rx6/iLLuQBs
vnOAvDwmIv2GdD7UZT7l7FKA5cTo+oigwiFKE1x9RiHZm8Z5hvMVyd2pc2hi8BNoTdAuuGnhsP9Y
3CpVQdOLnEdAdb3W3KQp5Q/VVMEZgwzPrjzYBJFGW7lZ3DMij+aumNcVEEap8Tj0cxVSPx/D4xPq
UftaESVmVWMJ0qyeOAEBoD+hq6WQcgPJHoMYjqXJLw81Iu8yuAp249AXY5Rj+H/Zw7moQL1dxxOt
jbvBWDWNCi5M7Yx+NomEGopKMo0PAEyQhcOpV1YsoGnhfEsgu0Sutqa642s1nIt6Xdu2nFgIs3dt
NkKAngavHxhF9lvSXLND+dLRlQWlytHAdXtYlBiVphkBXWPa5X+NPHEAE+qvaArcbMd8Qp/wZ7xz
fghbdaA7yOBNiber/qPhMLhh5DfVcl4pFXRAWTJpnDTPJu77ZhjtTfSMTM0X4smUcH/Yh/d1mo7H
5PwHrVMbIwp/PuQvvwDL+kI53iIBWhEIw5Ora+yux1xLgFUto/XADyR44cqDF16KE55U/P5ITraW
vRvu1xtSV+xNcnVgHy7K1wAH8LGXEaaBn1TdUWGWJbyTzkOUSLrwFPuZ2GahEnEZXtEu8U1v/wKj
a0huLxKavMroAMAjFYe8AYj8KSRZ2MOT/0FPlkZjWy2oeTxvg8AxeSME7Y73jJMpYZLp5G6G//Rd
NB9AEFJiGcTbIdinZ/W+RSh/I6gjz0Ap3vXmKwgkZ77Wz1/5jJNidEzaM38vjp15wkiDMUYHHa72
hqAZJmw3xDwWMERMvoUigcnYLAGZKnna55uhNdIz10cC00TnxNRHAtZZTBMCMhkiweETRcpLY/go
RvxaXG6L9zgmCglDYwW+HyFPKjVbuAXVMVieC+rzu5dhJ9KHr11LAK8C/b5l3AiyEoujmeJSWftS
H+PN/ceg2IDu9/XIce+bf3G1VZvLJ0f+/aWO0kZ24n8t2FaAJs81c7mDXrAZwlncjUrFg980mwTz
vAY4vpwocGHUhbJnNUPu1TVxAz1kVxMZTHW6rXYSUn9zJCUWUPJOxPdC1S9dfliLP40R3cTI6pDi
/7gXa6ZPA+CDZTEpDhyryTSot8bvv0bl4E0S5/Ck8P8lpTtmCuB83bncJnnDT/jjhERAArEa3I0b
fBG5S42P3WbR/RSYp3Dh+9n34jg3EzOh/xM7qy/vcCh0CB72U4kJ8P9XlZRX1qtB5y3VjZziBUdZ
BuCb38fM2VOQYltKFU1Yc9f23eEv4DsNUsr4QYe5Y5yammGpyEUWlLH91uvMHchRU8mBBI2QW8uX
t3u0Hq8A1e04qX30tvBfEred6YeusYbPAP4P+mOlcuTKj21xGMiQN9GgIhzVnpw9QHn/BkcNFh11
+JtysIO5LQ86KKyaakObuOHXAbhj8Aeod0ZxEIcnX1FWws9emItsDszQZlLmSHFs83cfXXiHJRDQ
FTV4AspjaRlDGPLOWAILcrjJfM/MnfGY/I5ijiFE7pJEpRZ4lGN5nedJrZgOr1g620HuZhijXZDJ
upQIpA2eWLqPmUzkdR4v0DUznrfSIsJKy0nwCF1mFUhmLqWb6TEGcZkzRgkTjlvOIco7Y+QAoQsg
4/fK0x0FJSevpsVRQFTs7Ta4XXPcYz6etp9gAxFA0umPTjrxG6cZhFLqo6qsrcoDxW7+sJvIlyVa
8j2WgWep2a2XvhMqv9N5xp4VGWdRYGi1NiTxHn8FKJgXjgDdT1fVAR/oX57hbfpkrBUbPfXypiLR
sDI0e/QxhKoo0GHhOk/lBRi4CKSDrDaFsKhiwIHq/NUQkkK30JpTnxmHX6rxGtKtppXMAY1nqni5
/ZibFc7sM9x+IgnaYd/MNyzzjX2BYfdVnBwV/EYIFfzPTNEW33bq2qhYpWBXOmaeRkuYWHHO0KUF
iC4q1mZW2uiYwQiQs70XupmAgIMxIIA5/Tl/HltgueSVhGVTkeTngLrPul16WWh3dxZVGDPZm34k
q1UvcNbiIsWhVajSDE2/7RINir09oQpAvSAgg77yvLGUHYnXkalUSp/hZrTmS/xv734I4rVGbqc1
N7Lsgc/xIMY5ooBlIAcXTxlfxkAVq6so4sts+pMBJmT8Gct8SZzZEHIXXcpV/g1jrvh1bgJHUaTn
zb8YZRk/eC4/IKGCysxHrK913ht0aGPeh0/BoVuV3B4ckX43Ef0TI5iRRo5wK3xZIqgrXZTfsvfe
bRXljIcohAbQ/vJ66YmsMT3sWnCrq4UNcyu6DLxKW3jFpn2p7SnTIGCVVYg7mJ2HU9lceD1ecDIK
oy5L3uU4pNH/mArHRZj/G092SesgUc3ufm65qhhSQYco4JWbFqboOh9cmp69YOitA/9UfzZ9WFQd
3WmZ3az3wG8PiN5seooqHpIhNz655aSt5LLWTfvdKa9byQAdYdFIe5bCo3IVlboWRX5IKex8akcV
jIbxLi+7HgXxfRNd/qMor7tY2/A8az0aBPO6kILtVlYfmAIAEC4RLqcSsw7lPd8wAzGfqcp0vhZE
6bfcPlx9GDV7D6/zzEkQiI/Js/KlYqhgY4HSeox7z4q45K1dXz8hseJfL7JlsqAwwu4jMWdbAatQ
CDKTCFKsE7ZYGGak1xzwj6o0wJx/jhR3m/Ou28EHzjjs7WgAUc5AxoxyKil0EuW/a+l6elOwqiFZ
Libr18HZUa/nymFDxD5aOFAZ4Q2pLpIL+8wuMEaluIdXCnXoPYhJRC6RIlVwYGmVpXTF46gpr1Il
Dr64Ffz0ucVyUDk9a+qZtsdnnRB8WEnLsWJovx4UeK1gCYq/+tB00CFNicB7EAO3MTGjdzrS18Rr
BLnz/dux7dbVgEzWcg6KO/RNFsKXas7h7k7xfb2MidQvKRIh/hH13eTlOZw22NJj2BWAvlBUej7d
dfHEo674kgT6u8p75m1Fw+iJzORVRyTSq12RujhD33OiJA30WDqdYjgyaz/zoEKWQZuZkuuxArO3
CLx5/R383Z+nUmDqOA1sRnkCSDDNyuYLDFpag8r72zEzLpbHbAgBUugYYTMWleglauHJpcubkREU
IEEJgFX8wfYg8Vj/DCxtuziakiWiBHFbpFNZY/QKP2Ds2bMaUJsby+fRgBYSud3WLcGM658ny9zk
+EuDy5ugWXlJs3jG5MQ3afjQ0yL38sD+3pgR4erTH9QtkAGllGsWu98c0CNw22xRBEJ7eEWe9rHo
bHuhwbN8/Tck23o8zNe4PlKgr5XnUX+VFbjkljhXFocSTKTrf1cHaqp1BY6w45WwSjvgygFdhj3K
wm2PKiA5a310Pz20hqRNJBeLXE5npAkz5ge5EhpktqR9kTM9N2M4SYtJ/8pRPxiEf9s3UooSRAnP
THGHoWf9TUY3FGAIBfU7Iu1dtQXoIebem2vJNXC83GGq3WzSrwqOfjgVj7vgGaKAErTWlsN20O0H
lfTUeL6U/ccjf7qUePhpLsczzl9luPaw6auABVUu4psPWBylwopkdLex7KBEv+0IE2dlT1Fryu4J
nMqJG9UwbSgNzLGAGykOkn/lw48GKxuaHSbD/axkyJTp/9O7RKfaxmonPn1UW9JFZuf+3xaTyPP0
nJxN0Z/eWWzk61XUti1lev/6eu3Bz/OMi5QUkJ+cNeVQoMXnACH2iixmaSc0j6ZEj7R1S0XuvqRz
EPajqV6MDcyf4vr69OJKJjt/f2M5nkiejHcZWEPVeJ7fJWHprJFFtOxBeOhdtTd4QH0/4Nr9cOCZ
0uUVadBC9o2YMyn9h9vv/3KSekZMbcJ/5NATwWBV5fgByr4nXxTvXrr76jnvMRYhh7xavnOtOd6q
5oj4/ppgsCUHeRxEb9i+ZXHCivF/o3cWYrr9D4yNyfd9iThHbM6E6pn3fw2UjKKL/K+i34GB8O0Q
KskaDM8k7SaL3mzQsgh6TBmpne9JzUJtpmUIfr+N3p9xeK2PpOXF63Vv93HGfEobenmRGC401cLr
VShjtbd8HmRoHSZBmNTKn3IH4LaIO4UobH0gOCkdhBXD/GUOYUaGtQ3yPKD1pQHldNLeBoCM3/w/
wi11rJIS1a2FehHuALWRLXFF2xMOOx4jrfNgCABgvNMyHB/tB5gZ90SSLBELtmkXA1tTLy52oYEW
QAE0WkfKXyeN6wLv8jaXlvVYt8fOObeqa5Ftw3/Vo0nwpgE6yPEykqgQa4ZQd063V0DebkruLTs2
T+ByYM9VSgun/ak7zDxJ++6Vh/tFTpInH2pITp1OXl/egQsrZ+Vqc0Iy70q4Ex1szQTCbE34tToH
da8iWnsBQAhmRbt+6hk0JC7Yzz+8qOu7qOedkUs9IATkULTAM+TMFmcdwvXxh5eUsIKXBPnxww0z
vEV71DE86kBeClRWOmFqn4kTDwFK3sxz2W8SgksKO5lDc2fsIDTvH6WjfpOqRQ7ukoamg7frecBd
K1NXNutDAekxRvthBcuv5759AB1ECasTe90q+WWqvpXpesleH8yVPwc2xOyIo5tiEAJBUaD02LOC
jLcXYjSdO5pv4EDCjg0FdTbb5Ny9onh6PL6FovCIHEODBa30p+GfUPYqY/evhPQ0HKKTWZTKkg1q
FtG3vFXcoIIeDVY/33yFm0ba3zRwSe4Vdw2ZZagSH+qlwyKvg49XQq10rj6cCVm2/shNhSefdJ4y
CyC3SaCYfv2m2eoSrbWpSN8z8BaVQcimJZTJ37yb0aJJYzPaLp5b2rcrA7I1kZ4Rt0wim44QBy5M
ZsyRWbfu848X3g7NnHEB1UwosvteukF5U1cU/dfx+BpOIRJKfQIV2VzCo2Tx+9it+HRkkAmoXTIU
yaPkshFf+8WxcD2H1n8lX0YLlaJwuTGiJCQ09p8hUmZKxeRY8i5yP3TZK3mcP+abm6t5rX08YS34
qNmKgiwX1ZPCK5NvtB3G5w4oYN5hWewzGJzPMzkpx0uSKuIrp7lWIZW7wUaYKrEM+V4dVUjvoaIF
yrYC7HXJFEI7+DmynwMyLmeSsgyXUAQ7DdjWPG4HtC7kc0i8aM1NiCz7zmIb02zJYKATHjFSqset
l/YL3iSQcVAjj6F3z9a56LGiQOmueETIshaAON+oh4PNgXrnEUTzgnmet4q86zg+62yu+W2xRKVj
g+wOcjAHtf+KE6ijvjMwklMaVHxzb+XfnCebteUk4uipLSW/tvaO2o/hOvMEyCAfgB/fbriFZp6g
C9udHLUb43CEf82ryiKgJInLOryio6K9+yl3c0d33C0zuncWv23hnvpgQ+d+ZnbHGT4fKgoonhsg
R9twLoRC24naaaiapbI0g85ODHH6hZyn4Pq84vamkwhmeLF4JPDCft3/HmqThSL8tzmopIZ9GsuU
KKal86qMDONZWpRO1tCPZ7hsc2zWQxhXHY+2HhcJbkbEUrWRfZcGMakSWkeEO/UAv5A04CgnPycH
Al1yv34R+WEsiY2CI/4jMis2M2BWkJAchbWWIEhy2yrnPUs6mP+7iegnucA7kVtAUk7Qbbv7+xEZ
M2/hAsR4ckgSytYEKQYB+ctTa1p52k9oJ6zOPCjE55/ZaEEH+8WbZY5OOkyhFeI+y42UDbVm+ZZf
1P5o5Lik23tMJa04l1qgriAXRVZW5bOhMIPZZNDO238nPdwatw6hVhZh21A3Rp2ks+I/T5tcKKSd
DYr9P9VQ1X/j9p4YvMUovkb9Cc3ESeA4oveEHiH9ywmWGILnzoggbbbLX0gTUVt4as8hx8DkPYJ/
kIVBqm5APK9doYldp7pNDlaTQhTFRkGOY1b4YPiAZVoDDdO6EKy9Z6Q6L7mAfrSeOrLapBAlwfwI
SjW3/OdiOfw/FbvziIN4NBNwOmJqKdxNJXRCnJPyYBb30Vw14aVzpJQubTaFeVDWM248MzmEZVbQ
ocMkWG8R8ipvqaar5/ly3NELNSrOGRzBcp4pIx/kmE1zl5ecmENaCKrl0du/LWdmMh7XyYfQHH4r
uHFFLAxdDuV8xhut3GtUhjl775P1CgOqwNYOg3dSau1J2NZQSjcd8DlDFhfrpycnMBo8cRaYJ8mB
XU9aRz0+AMvdWbCfeqPiz7PSqcWbs2I3HHUT0JfaiJwKIHC1WguJMBpTVvrJMvlrzS9nCZBw6FZS
xM4dUGQCq1dWvcaReEhHVT8G5DJxTrugkbeuDQpBiNArGT7q36BddCZU621RRWc+zfzXujMvdhVD
fuAKuIPvX0Ra4JEji9yfBud0DN0Zv6C4Mr9IQY+KlURA7RTIzy15E4X0TLwDiz/k4gOBirsJLSzb
JdwXDRkDBmkpgQEwT8HXbETovD0C2SktyYA3fJFrOdDzRntlAdpnUZxe7Z0P9QOLwq23nSsUrzTO
kdxpvsp1nF5HYmkTSgA7Cu+beFJq3j8g78EGddUXVwavBU3//AmNpeDifYEeLt+USbPohruLUgbJ
U9UM/0TBzD6gOvLWqGBfnZYWF9+lauFa6vBVgPlZiieITeRJVzgiBrkDlweuSU3EC/VZWl4ePGt+
y/0fNx0qYgB2l9GPdjmRXksIoVOAKiEp4Rby8L+UvQUUjugvIvsuzKe49ribix+CXS5ryrbQmfcK
zqlMxAiJ2pYlA60jALP46+XutYvYLNQsgnxDkife2i0d+cnW/HGX9A0pYCCEbGyTr6TLjnGq8mlb
WWDpYi1b0jHqwSxSq8KUXpeSoZKLntv0JNfJeUsoQHSLVTNykJmOYQHVoME/wc9fUMad1BpfSdx3
Uw9gRcCjzMVLruUyTAlnUDShQXG3vf13jtTRsIJw183HP8KjzMyLmEby6l3JQO+R0/zjhz0FjeAZ
fzwyRh0VTK/9V8/UmT7vr8O6RDfwp4BORuf3hNQAxJZ0nb0RZ1wPx/YqXnJhRn0X4PZ9Fyn0R29w
vqNWBpW+QfahjDWE11h+VL5lZdG0ipWiZLP0XCfOz5lymHkDTAmMfqEny9KwBZ6TNNpdhm3XFOQH
kaosXVOgRXUUjkOaIC7/N10vkgYz1bSNfnsDxXrgrm0Cj4lszoor3xO23zEmIt8tUAaKpD39pAMV
gW372JRrHF9lkkqL0atrfIJowLWPZWnkb3Wl6/PxUkRK5f3/1PWhsKAlX45HMu3Op2MWaYMvT0yE
2kapiqUjpAZENdPVPQuxtEwqpGEaLl7VJ2k/wEhhPS7W6w5voHNCwSjteNnk+b9LvPYXMt8Qr9q0
Sp+6Iqt0/MqHCGVlL92f6KSIKfkE4KJB6NdyaCu+FvZ1eryD4frxpAzFG3DgIexpP8+fhRSgmmmL
pMnFvJABSMVt2rSll4pNy0yo/0Ume+JSKPYBLa6D7qcGu8M6hXIRUUQtAqLI+cJGVNrmpamo+p6u
nLyRW1kFELZb8QO8sEZvfXgZi7gstKSvThqD1fRhy9VZo00O9+4Gfds6huU51v6aCwBbN1y/KAox
5WO+pe9G2uBVw4jBIayuXK5ZvgBaVGYi/Ct7ov5mh3I5KMARC1FJ/FtSUARIxkgr3AaXrU39B4yQ
EGJ+dhOnp2XC5+a3nT3Uysbm6WTKpwfeZbpLGbmcU2o6KEOE4hntdm/syf3YM/LQmEOfsWLgFszS
GM0WX/QMxg52dZpZ8BQactFXFLYIxsOUp97d+mYhpgD9oVltVpeoXgVnenw4Yx2xycHMyk9hc9BF
sPQLGEN+sZ3NdXtaCZMQwCblAHEFA5LG41cheSpFYhHeXOlSccRQqEvioMtJJ2vcVZsqVTJ6gqr7
NDnOM4O4UJRO/uo5ViIuhIdBFXsA3/DuK3jvLmCYSlnnc20TFC70e8q1V8vQZBaNf57otGK9hPFP
c0k3NrqftVK7SgbkdMZjd2fJKzZ3/jl6DCLGsUd3r/1aKaKzuA0+F1UQHaax6IEpfFppE+CqhUD1
HBiXcoW5WftvhXA4vQfiUfBvkfBWNFsbbsoe75Xu2J4i/TXj3/dyV6hHt2FL2a4NZnTSaerVFcKM
SkSbEDXw1Z4I68Lx7YV4zbCHnfmVWtC+l1boXAUCbWGDTOc6w9wLGdMCgTctrPPMgIBEzCkVKZg2
7abuRcS/p0hZDLvaspBbo5WyljKbHKNARYbAzkfTHuwXZbuy82XKNTgBRUMMj8L+6LLowfrx+HDo
2iphSNpkP8504Ef19lOmaN3MfRa0ST+Z8JhTc2hW1hEVgs9HacpTJ6CC4DdtIyr8XwncypK4zC0D
KUjOrNtuNHg1ktSmalmkQkgaIVw6mXb7P6Ua2RfW9p9q/gutkc4Vd0vpSPPvJ2h09Vwjc2hKenkI
SgzrqixAx80ZAjAZiaVNGaQ54wkrs1OvxMf4R3XbFQpM8voQStsBS8FsLRTk2SBDZhmxJ550hopB
HIwaKE2ZZ+/DlNbCqld1BH4kEgr5jzNRwj1WKzn8u2vtI4I1wKPZHhOix8Fl6n2f6INSQzcT0c/i
KEeFrWaCe1MMDcHAYha+sEuIFXfKsVQh4tZoXMuUg/Fw/nwX46NvKc7BRVexEw3DXLhzlU9nwC4w
idQXyBzc9xyXGzH1Y2dzSqU7qLqZ3S0sQ1G6wVQ1HhJz/SfBsYSvuit3sEVm4cbFTakQAb0/rnQ0
cSGj6DGtrtnqJP97n9vrOrGoMPq7sheN7fUJ0k1l6XlS5fFs15VMj0D21Vng58bNHRy3oeL5V9YS
Yt3rwkkjPoY6y49Orso7DkSd692hlpbKJYoNGKw2aOxdlsq9r0GUXuk4ijHDyFd7Y6z7wlpuPoq6
fYqMSxjp/SCwHc7LDjlY/5/ofEXvOYTRBMcHol8Wk+WZIFsxn/Kyktmp35hmaQmp+xuiWtneexiG
nyXw1RkMCy+CaDMPVARAjFkR3U2LNCdvkET4MUDNMqrpcny3+pfrhcckk5F2Ed8CsJMwxnUgEe+K
k9bFCzITIhpKRtTA3f8Dzn5IjyUEkhprLI+CyQvvE7tTo/h1JwK3EQSwn1ypbT9FubKqV5tIi99I
PzsY2mLHoaIqMi3c9kZdLiF8yn5Uu0LRdmIvTXK5Hv5jMmDbu3YbJde3Wc6BGyPTRNBtgcfrnY/D
J1c9xM/3JnOoOXloRcYbxfeMTnzQGWw/splg7rJoqXDdxJhG1Oe+KD2NGWuYJNJ3LDwcHHbBIdMD
tzzHbiu5jxV3NAq5xyVKRWM/WOLNz2SdcpUJHPmSIR833U2Tx5ysqChypPh9hsYqThqgsAlRgjFg
U2+MF0xDo87gp1gRgDE+sYBEc5yuhspyCz/jXB832z0N1z9T2XAWixXR9zgj2mHDjqrDYQZWdytD
l6WrPYOHr9XgdDIypshTzihr87v3hULg4g7U2gX5fq+IHgBqy2eh+X47M9rBSkug/lv5lASZ9FWv
qUrYpREd01xaLf4JoQxQWFp5OWGOevG7Dbxt8M9hOUMGbdWRFSwKbePvtNe+QXrWKtRrxAH3PnjZ
/2HO/airBP3U2Lppx+dL3VU+M8XSviJOCFsoKhwOA3t01YsyYRZ35AKVjdt7P1G0+PH4JzdfrSNg
t3yhEwL5JbtXtpKfq7HbbDdcizAGnhyq/WA7JYmP0fvKYDwqB6fmq4rIdib01wAk0qqh0NFnu8LE
4biIATlalvSYnZZebcpmfw5fYlLnDqgBTyeUsDmkNpEezQC3ZXYCL8VQIAazVKb5VwuxMg3TaoEr
I3Is5Uyup/9MpDNtQJWMNQf8IosaPmSbjtofsyqx+PUHaW8DATDI+liRCfn4G+5tbbz7uryyUojs
wUpoR563vh+7fQjz1uT9WgFAOpuPOO4XeVxo6RglWMx+IakkesR+4OXr6DSCyHeEDeyT8WLZXdsZ
9qlF/aBZ1JYQeDakIDg18g3gshV/B8UuyeUNnQ8AaEjXv8T5JUjlZzAKJ9kCx86qfwgPHBsnVkbJ
BenZ03SevFoX7XuTr2KKJ/7hNv/NOrDz3hCOM8c6u4MtraFnFDrOgIAbaNQW3wHE53om0eCullCa
N0G4GfaS7e3nzo8rWggA4wK+bGrJZbEVA/rRrfSSiPsBUL7QhzyZSO3gDXFLz6qJGLQqojqlTkOp
yNNGLQL5ugFhHUcQzY2T12nn2UX/htcplAhh3DiDxYrRSvhoj/2OmmUZVJEQsA3BfhFCecwsxF+r
TzHNVY9gHOyzY7VxPUTDAVwgkp5jbgvbalYaB44/NZTB2/bS4qp33DoKpQtVHM35J+3gCmvJqnRR
hLd2xQyB15HTA5fOUNsYq2cwXH9h7LZ8eXx+FXnyI6cJwPZHncQsZX5SmiO2kjk30WBCOwYEwk7d
KoHOTLPPlavhHsiKpGCdKD4stZPx3o+uySLxItFmTle6uGiSDWunaC2mlaaclTNdRm1L/f4y2j0n
ilRjSrd+KoEcRt9eb3XSc2+PJfm8ggpkC3cq4mTGBWSqlGlULV8Z332LqVlusEHhvxngS1jJoboi
letBVJP+OcZNxl6Oyzq0QfEm3csqRtXvZVxbisJiMVO5aDap6lIOyVA43RvyBgdbDCIrj9Nld+jR
jVLHuG/4SP8Nqk5Fv8F0hOvVeMitPbSlYWrBYe/jJYeWtu1yHdqOXpcjltaQXoDM/28hiAEohsKL
zngwuw1nXWCp6fGaqsw6zBqeLcqgZQb/FDdmgZ51YcdrMEEzfRdZk4mxlDyJGppv+ivCz+pbloBE
Ypir2b2Jjc/udfwMgIKJOvyw4F/p772NMQj3x0n9ZX8HatoV3YPq5eopuNmxDxlcMflo4qWXYpuZ
qWM2I+kOERVvfyg6HKMZJHJYQ4dSpD+gwEGlLvpRcehGabaZHq+beZ+QDdZ8Qp0h0i4uAe2ttaSZ
kvrc6TfsvI8xRsg46kXKiPNvREjbrC5yPoZACOl7yGKsS0zMwMKu6HAzvp10k0BeK9Lnutp/8nWF
G8zUho1dmyJcxPQp2+i3Hm4wXCTnstqs4qP4xSSk1yuMabZtA0nre7EB1Mjf3wc6aTP4sabP8Um+
NJXouBZtcI7vMg8EDCnfe5SBLy2YypMh/9OaJmzlIanbOEAp8jAZ+e2OUfYwNxV9EodiguuHFGNw
BuvyB1URpz0rnDaXAa35Bk7oxPk8D5VkrV9Gankj1zyfWSobBFZEaYpSAriEIivjUWKH0181GY6G
nxYzBO7fdB8j4djmwYQpga+fnsrjVD5qsT2Zi4tI4mCIux70l4xq6lNOaHINSpy39fNNZAUiNUyy
QWlu42pbg/5ApiiNdAIiJWkMgIXwCc/+dcxmHYEgp3n4VL3/7/glDfYj5/I9GdxorIfpbD0B2ho7
vhR/TlFKNOkSXb6meL68AR8sY9hZYO3biHW/KWGRHcJmmQfpY4mhK/ymZTOISCQP/2mklZZ18B+d
BhwgvwH+YbxDcD8KYp9EeeQMqvNarcG+Cgxx3w8akmDQsJTfLDXHlzP5YT5Vt8mDy1gvvAd4KlZa
n4DG+o7q3rGyiZqMGQ5z/aXguPc+djwl6dlqGH4l9bXbS18AXMsKoKnOwWvRsF8+XSL1amSWSHnj
MfaSP7hlaVvLngcSKlQrAyFS3N87VR3oWUTQqyJZ3i8ngqNbdF4iws+yvirsXil+m910rAplO7Gf
N7r8FmWJglF0FynOIoP7+/xdUFEL5dIhsRB4NScOxRmfzdLKQwA5buxOm4axYyaKPqAZLlDjzkGP
HGFpsxWXwB3I+nl558H5olf3CuBG97/PVJ1Smn5nDwq9eDXtu5toKWNz56uxLCqvX/XUxC/6P+g8
V1gK5Au6HqzzEbntnEWtQNcETtjlX/B+Hj0DaGDHKIy8FqSwH7CUQczZyvkAmskNimrcpq9uBe88
wSpqXxXUqCJqcvX8n3AR3iayMDxitmkFTxeIMlDLWCvzhBk4XZLAxkkgKPwNSHo2fST9rSxyA2cS
V3XgfDizOsjgB/Unas8F4vx9JlgMwMpOaXJ+tdM/xlOAUe2f6FMB/zzSehdK1Fm7t7iHuwjY39eN
QnF0IUG/ndrAHypTA65tzoMhnk5oej2FBz03YD6nNUhcYJSjZ9cND+2wHr2XPFmS5ueg1JCsA1wt
b3u2Xbu5kGP0Nr2q7yG+WQQa2CrFaP/7HOoXmsrG4I8WQ4TlU4r9+N4cnKrhwp2R4pDzQvrAjotM
LRNaoqtSh0ajEfUa3heI0E2XkqUDuYJ/BzAHPPrKVI3PSG2yfOQzYt6cun0JayBs26zr63U2eDuX
K9Vv5WQXqowJCo7hFPF6ZnpypcHM6EuOnhe5/O03+IMjf7n4OfI/Jzo5QcYSb4PdGzu8/pYTLtCf
G1SRkJqBCONbncLOxzPqmZDi6xDNF9ZBsw/MzqnjQG3yohZPo0dC+iZrPSAbbDm/KRyvQ6mBmrBn
iqxyUfmBrn4E/D0NUhFmGC1uKUCLQC6Nm/Q3PU3COozFK6pwla6MzTMxC3JBd1d69bhJzEvpIjo6
dK89P9QwfT/APJqnvcmxlHPK3qBgQCDisfE0dnhXQu/uhrhxffKjFsHW66FX/uLE3j2n1OQy64lw
tGxP/3oktWf2rT+uBshXbfdts7sXJ25uEcmctEevSDnwmoN/6PQHef+KmSEH81gqrD0Cim4glzRE
i4Xr4HPKhm2KnJaEodsnXAa8Kv1SKmqAaHZROPqWHUyl+MIYlujEDYX8xLJjPcE76DENy390N3dq
lbR/4xDobBibKI2ega47e2jJsi70Wo0unGdgzPbBRj6CBB0GZNxlQ9yHOf0353X4RyBCqwujKGqE
Wl/yQNHFKDtA6QzzayooA9qL6eHDdenTuW9UwjvG/n1C1QbqMqr0sHexGPjKqNAIZRrnyuvwJPko
RAOBgV2yujNwU96tgKdUqi6AeXxceauFPTR76a1K+XuNTLo0R9mxeHFP2MfWtOllBupFpxAbQE4l
gibRA/JnJqFV8CsvwVqoqZ403oAG0eoDS7QTW9vP4SvL5YtgADh+tMb6N59IIvj6Rx1lEMbDP/BL
LTAODoQ+vM+bO4MUPKKsBTaLVAcVustmdt1CrdY6KtFwVI4zYDB6YSrocMTVDQjnvc5vhcWW7ee3
pKA8pVaGI5cZ1OnMGPagvp04y8FXudu4iRaKNRomEV2XCfbCaX9pthMKdEV7Xlch3UyAzuAMq7A+
115OrrDQN/RLGVhAj32OQAYNhkx85QJfjhaK+KUcxqQaPMhYpUy9cwDqAb3PRWLALzYXo8xTwmRg
y4OMUWCWUgfkqVW0rbtAbRgyqWk1H+dm+6L5FMTsj77Idci32CqaZfwRd9zfdftKNMJDExIL3ncZ
BZ51YskLjBp0PawOyKX7arMoH6KOXDyEPQFTpQmX8DgsYHPV24fBahcAppLNp+s070gSv5+pvFyg
tPCVOADquHXlPwayuu5TZ7Fg/Lrty9F0X/VcD0vTRCJr+o5sdhkPozvRrmMkiGhHSkpq3G7KCMzz
Mw/7VmX+WcGHKM9YGLro7FzJgn/Wy5gGlp+FvJ4GpuEwpA+nt3TQGWhrS3qrxWPGi8ejjMw3vy/B
DDMSNRUuEhjQlIAgRe7ehvDi8o10ZZcxDAMQrTVEwpRNcpiivQ1T7jm5xYTaXvDskzzb+QBC9Qh4
LUUia0A/i1BO6HPJNUnl8uJuKqiwipVWs1HQR69uGKW/lC+pupggYffx56U7D3oMXEHGapv26epk
/WwfBLaTPM4m2UHFIxTyy0J0kjt4XY0W13Q1YwuGSPPi2ggpskX2MYBS/+LUXscP97rvU2KHXeMj
Od1sL1LQiRDUdudBfdcUwm+13AAAkOLsKBM707kxSo7Yqaxqfwuo6hEEMFseNWfEmIYVl7Qx9u2o
gY4MpkCRvonqZjI3sTWhsiXpIcXqEtghXGJKc1smCRARg0QQxV5YXxL9lLRwyslwyCkJtUNcF1YX
nq9VFKieIx0Kn6JahqabFhWzdob0Tqdm1eEStSLDw2DLu5W2OlImjB1iffN1Sf9uvih9fOl4EnqK
DRN5D18Xzt+DmEFDopC6eJBbK96SfcZjt6M+VzFfiIrN3M1Fa/z6SAppiGwZ+bEQ0M6YqCcYP+qn
WensaZbxCwbRDKwTghRLJiRPWcQRllXzD/28TPUHUhpatqlwUhVCZmuWY0NZ77DLIDUiLPzW4H/x
xAGSZFQpsD+/n9NZW0ClEsnMt7EVfZcLmmCNoMeZDdIS2V0H3v6Wfsx5uvEdz7c9QmpNKKFeJ+g7
pvs4+4b5FrWBP9/rWhGJOXgmjSjdrDUY3+DzslRiHux/yCS96cTFNmhYwijuUeVb7ecPl6ZU2GNq
wahcPeMh2bLGY9Lv7eKrEz7Ri/IUUpRme8APn7M5ifdRO9OilAMAaUZLuxywepPyUBT5rEYnHeGU
kS2nXBXPwbxCc9pchaNtSOEa0uZc0Hk6WSt2ySdi+CLogKMgTPwemliFC9phVcq9SUJO6x0S7r2H
CUGIBoI3kBbHEujyektZF5VeHCgFizmFKxwqPZzT2UEiDlBtx0eDSq4PXsd1befGWcLg+PuSjYq+
VrGw9tKuHK9g29UrYBWc8Tufhv/z5dzXNIzVdvE4L7fI3UHXBBv3BbQT/N0127BoaKn0efL78kGE
uJAXvEzla5rr0m/VcDqcHglimbqe1U8olLTu9Y6KLJNWZZj6NC1qeWLXBI/gqyMA2dIqjXEg2mid
KxZ6M3dhRiedBfV0tWlCL7eK2YNIT4jh+ItaBXFq1mzaWKcMKVuom3MhhXGDvGJN9kKA0vrsO1QD
srE+kIqtVoVejTPs0yx+33P0yE7qudXjxKDOUSDMueaS1jfp9OkUEucCcIWIC+Oo6q2DqfU5AHNS
2jdo0fnGi1b7c4rsTa2Vwy9wzH2G0lOo4s+nyqrTeoA9r9MIz/Jyfonu1fUpAZ682HVwrCQvANQW
FiiwoAag9MLEMBMmEg6AUOS2YQk/nbOBuHJI4zuj64PAyDBXAUG2QgK3o11agrl2Xn3FCCsvjiIj
t9Bkkom3tPuwzTKjTuf/d+CA0+Y6LnQNrXl26vnlxZo49rKvnxUHOSxOQmaDB7kA9xUdT8l6rqnB
XvFYjaipoLmKfQtRk8/EBxJjC45x2aLTnDPao6W5aL8ssv4mWlNacYU969wZ47UiGv4AYCM5JyX+
bqqT8bGITeWj+9F/2FbPgBGVk2JGG3uwpg3MUuRsOglIzZoZ3V4X3pawYblXhq/tJ9n4EMgMprNt
YHNY8BHk36mQ39mVAKi/NuMa0R3WNH2MXTVTREEnHyhH0ESP49QJd4V88PtR4/5XHIaCYbf8ZNpo
1gpx9TgBgU5ZS/dCSzk6AMe6amHuH3DVPp+QNyJiAkHA6lZ70Hogn8cwZ8FKZcbrfolQVAjsECSa
jJHJVIm7/veQhGQ/rRPiTLXO90xeVzpFaP0RN4C4e61M+kQHHSEreMcI6bLKsDHYk+K6IXKch5Lt
MBaMEouNrwJ5LWgcBGzzZNpmNI4YtbejqkQsTBIohWPArsEC+BZrefIaJsbIiMCo6W3HeiDKPAGA
1wJb4RAODNN5na/MYOAyWYTwlK7XNzYLV3JvjDKofVVK7G3rXFj++5S74bnVKN3v3zfYeV16hk0c
P6vmgf02IjYslG1yAFrv04BEz5LMvArk9iN6GzAJNOJvRQn7WpxvkJbVDEDand/8KP356rmqc7AO
Qtaki1PF3xyrSCLp4VIzsIdEj+AqEcesUvb3Nr9eeH99PHEdwuruqBbiz0vePUG7u/jh+cleZY0I
pF6qgnOrnJdlMVtMTahSplofpeVlzsSwUwqOVA3siYUzmWYeM4baOmpIM0trYNz7O7388anerw+5
/2j5IPoq/O92WmCguPnyVLtjP6XyUmXRM8BGq38j6ojVk5Iof4c4cC385h0b5a6wuIdf8ZJjKX7e
gHypOl+cbcTeYMa5YgsQlIqREKU0I6IvxB5jBgYGpH99XwV+G5VL11LvKgLM6lIwe+dPZ41aZLfr
y8DzDkk3L6nQ1Qhfjy/BOYSNHmBTfsUeseSae0wVZMrkIX4+PBLqtHOt+JGh5V2JFUb7HeuZhO+s
qzPUVPCBMYONmRuifGRS41p7ewTMt1pmMKQpJI65un0ZIMyZtavfq9Rk6dd0dyHlm/V6naPg+AMB
tnhcwtXosdbULF/zR1miG0tB7hlfG8pFAM4E8T8eFgLP1p3nNMArYQ/jos5oKPjl7AcUa758cA9r
onjCGu/ixDBno/ssdIRIHDTvtjFMA4cX5kwMrolzAFEh3OVILStJBA+FwC6hRhTLhgyMRvgX70RO
jDs70t4cSUFfUbVMuNLdFLOev769e/sggCSeNW+ys0FvQ6JKXomZM61xtfgTELmZ9yPlF4J0BiOl
HZy/GNzx+bjoY5MvAR2yHiry2QHGWmeI0YInKZ4s+uVXapCoohi5kcen3x2TOqiCP/tqksc+qj4C
y2vp6ms7R2eOzLRUAFqv0i2JYZtAOnndfAdUTTqxdx5e6BsyYdEp7dWZ1AaRUCprN59pPI4ua45Z
dAVnVPvoiIszR4MnnGaxs6cqVnVZkrjeLfl7RLsdwlR2uo8th/QelKe4wbBExh4jL+kXcAX1V9sw
KFT6JPu7zowaLcyW5wLtdlyu1qyZMHlbtI3TmFPlhc6xbqAt424JX6ezYiOoioSQ2hMEZHzZorOo
dcEE1HKU16xdQUnI5lpI0imC/upgYtKqgOFxXZx/hrzV6jHukokqrSbr/jz6o/BjY9uh9HAyitFs
nR7R3S6SzFLJyKknhHg8FBBlPcSNKcdfaIksuJ2FtmEX6ASPn4yrdOK0c+Q/bj4G9OMmif6e1FyW
Ay8ypRbkj1GISCRwrCd5VycDogGQAq6Lyq4MphSCiGoB6gIRfWK9sEKAF290QaTkiOv739fniijD
iOOUMpYaHVeFVbUN2nc7rhZjoDneWdUMfF4ytd/4Jgl/Lfnkm/KIW7y0zMFsMFDKIijy0cYoAHJN
lTZSgf4OtvvHnJ+7g869fXZmo1+u2Zz8ISvhtg84MG1FRzrsFqBxQ6pCQGMrRw51WxwCmuH4Ow+P
8j9ZwYQZ70PjNrjPpwyMVvi0ZG0zvtR02L0ZQt7mxBSd1UroKDdOzLhMvRc7a1dSIF+P4DRQhzvJ
/xiNX73d/FWPm65/lDZIdeGRqdnOZiF55Evoh5k0bpZiIufVtdzwGVhR8BfUmvOWUSyudF5EWkyn
GYM63Bte4RVuEtWXx3RiADrb3xRl0m3q3CA7UHQzyWMObbZLQdAsPza09v6USkamadTGLOvO7pcS
o9PeryIJDtERhx/uCCgMx7NdHw9bDgsgaoifYFctahXQ0o+AZQH5NTsNWISfdoDL9XUpcbp1ni5L
UqK4hhGK2Yw6V6ae+QyBACZriTfK8DlfhkF1359DtXisQ2ZeXgcPJcJfCg9oKNcX0yWZZMXpPCeW
V+3RTitft4lRJHRYduaX2uOgzSQOPgFXkAyH71s/58ScHJWbw2cu6HDJOpNhJxF167yY/sZSbw2L
wCHxDyLH2LZsa3i65QoGn54MfIfRWX1JIvbVIzOpATnT6sXZDSOiEMkb4eQ/SxuuC16duR/lHG8s
0pyO2kqyNniltL9EGCHmgMeQq49Ll2S9MYNErz1J2J/SYoThkTpfFx/8+CMLb58SuTVw3VfK5OpM
jAssOoqIUW5DUVijAxdkKVQ3hp50cE9CLQ490fFVbIaO97sQalo8oty1butfPq/Xbq+rASIy3jTW
9Gqfr2xbscEDFNqC+Nt8qvaCdbulNRLt+/Jnq68WeAKLySqcEuCw3x7xVj2M9eP+5vgZLmvaMeJE
054kWC6WpbWtS2VUaoQ3D29VGPL4eGKSTU/6NOzAGAJbmd7MfPF9CmrcbfZlItjAbezpKN4r5y+G
e2n61qivDQaTwn4VBxvxBZYPfvGit86f4qcZA5ACpniub7n7CNSajf4EtgltekwgC6EXkvsuY4lw
QHRCNpULas/ccjmuLvBCkMR2xWK7DI7eCpVqdflfxcvlWRB8KYKqSuSMbsx2f7H4IwH+SL/rZY5Y
9PAk/50es9Bo7egDkzq8L7340ObsBl/4Haq4OeimGTvaxn573sjlXvgRnd270EuHI3pSlKFRRNEy
Gj9MBfqi5J23T2GNeqZbsLdNitUgFtGWfnuesuCzaPnizRwVOmNOcCbB0iTfMp/mLBaEvSPOvPkN
aT43gvbqjaw3TG9m5hbw0L4oSKeqiSgOB9DBXl/36Lwx14rXwNRkhk6V25xUndn2VBRpOvLERjb2
snZ/qfGlhZ8uQK6pu2wRk8jLEamDs1Mi4BjKXhaO8UWYxfqBaNHXyvZ5tR2MT4r1UD4uDD2/0yXx
6gfNsqYZ7sQ0wyDBtEcSDkkYQ/4wBFVi/CHtPZkB+y7S2M+9QQ7zeIF7Ez3FIAlMn0lkYV7YFmsU
5Z+JhKMNxPD+TmpKkm83yrUTjn0UYMuNkYr0rgPTWXkSPf7nsNKN9LonLEXG8dEmu0+vKXvLeXwF
B2oMDjMMw9c4x196BvLRKZt5GfVXxzwZpnONrcfpL7LSVHflYyKm/bvywJmItqXRyjbNmmS5MMB4
iOFD7Fl1IQyQs0af1OzIFGXM4DhtsNc8WO+Edkiamh60RJ2zmdC+LePa2FMXwe8n5FlFILdSYOD7
nN5SPqD846avdcLWTIXVR03dIq1/gAaREU2lyCETnFXC7HpeLjS7wc3ogF4h8cDZVNxClS8zguJ6
B20CRLs1iG+QUkMFAbCAC9AyvxYuqoOsHJaEKYsYnBsceOZXVP67n/alhZAt09btxNpz978UuiCj
x7cvP3yyKvkyvfOpapL8ypkaCgyVONr8wd0vaJUHWjHPRBo6l2obEH3VoxAtDptAIMGj8FlpqVfW
7qGmfn2LGntouRNNFDtxbpenySIfPCgCB1xb/vBa0aLrxA0YdQWQhMVJPc1XrJMiul7txdFkpyHE
RTWW88KIwUz6CBh+iuLqU9aDJMcmgW0cHkKFIZSrZGgRTCGd8kOA/dygMyFQnsVhUlQWO9i3s81A
nNnm8TgXuONhurPN8AO3fy21sKP3fRRW3Zt8fNV7694BdSJZqXyOerh+ofiuzU1BBXLMxAQ6hiUv
2HCC0KkRb0Sk9YFYUkai5sptYHra0qWymMUz+M05aQZ5WDEt5X5weSEVJJKjeo5RSjmYadWM3Grt
dQJatoEZxB8qXkE9YtvOZDwdaXwyaJxhUuPh1iUAs9WBnNAIE6BWugk+AWuxSz3WEcPCeRgzaQP+
CRwrOipfKS2Qw/YDkoaUP/lLM1ooVsWWUzVWh/8xSd5/6Sd8AchZLfiEJWOtcz+YahKv850rLz4q
tqkmR1cl5A8Me1J8U/+KQJW3Mv3Mi9BUCXsj1yiBClXn2Wkj87x7sUVBM75z+TEfGihqIA7JN7a5
sdcLrJgl5tqM+Kh62YaKQwwLXX93ykwnepYNuBukVBlnpEK3RDipPgcHQxrX6ZLHcrimNAyaw3DF
pm6W9RpwNKfWJUmHxtaZMfNGHisdUeqRaL2QGQ2EQ4S/4peozX80lRBRHtTjHM+ewLyQ2+AEzGB5
9vJZjmzplnLn28ssNk9fD0PNWqR8gbwsshxuN9ZpRRkeBCQsViJC3YSBVe60JLhhLQyM3gTGL0ns
AlS1hkaLo93YQbnjXPNafe3h8Y5yLtX7RR6+bcPcCwsQM53VAIp7Ba7WEkBxl7ZK5tNaQWFFoMim
hPoXvnC1ejRpgYvmu/RJpHTN7nouXf8SuOk+b1unLcntEVTPHEibfF7lx8XkuMfG0X8J7+KADtSi
ZAaoCZp3MhZYzTAIVaJOPBWrwe1Ef3mgAqemv8nw6W504d4CXtd64O6So1IW5Y44Y86BNcaRyn5q
hDbs89X5D03zaPGNzt/GM6uSufqyHmLGdz1c3/yxr2JLOJDjL4fNmqRW91TmhugydGoTBhqRN1F/
S9bmE6QR79cmhZm3VwfCibPOGavQnVzdj/8xDJ6F7WZajLNWWuiPEGfaq4EDNUa7CZCuW1IH70oT
+d5QEWmqB84fH1cGZqra1Yq5zKcSJogfuMqbNGkzlHL75vzNZu05M9eV2KG1/ZsxY49ELAhVpbT4
B8kVRsp8MzCKoPmKFAmOONZO2bPtL5jCg0ONpObpr8vNcoXdo2sivbfNNBNj2DGeIls7pZ9MxWpq
N7DibRE6PKes/lKeixLyz2b1rzWq69Im10rCoBDpVeYQ6gtyDNTBU9z98Jin1SbLWCWro+ISDcvB
JqGuEPKvOKbnDcwIh2SQzIWBaSDqFBR7bdi41VADFpnEUKUfzmAp4T9EH+dET7LEbzjiZYCZz65F
TIipeebuQ52KX5Nuth/2DFrBETTjLFSnCQW/23Izw1wozK8ul7GdVudhjR4HyA9fT/tZrBRVRssl
03nKLZKNJj5CDkT2cJX1Th63Kqg515WtMNlbS5yQQUvZ9Q+oil90UZP79Vcxhxjq7x1rWSuyBLN6
GJLhPfhP2Cgzw5FDjOoTW/x5VcJZg2yU725TW0JbMd+q4x/0FzHfvlQ0ffdbzfERCxc5uKm2WmJL
DknH6NwL2cuVrLD36gkGAbeCDJKbLgje1jPsYq0qb0J7H1qW+WnPeIHsMJrwPz30Noa7AzfF1DPM
Yj/ajzuMgFW8e5lXQmiblY5U/TiCEQF5JK8J84lzbs01jrBvIY+h24nuceAHty9iCkg1hyFvkGzY
HLgVi0ltSIy6VWgLJlRw47VnnbD2u8CSdMowvXRgz8EfYiG38pxSs0vvzjjLPhoiXqtsomVyE2DA
Mzfi/uv5Du/mptl0bJsgQbhkZkWzP9e4+SobTKZ7cQ7ijUpvIqNjJWHUjlnnOWgakx1s/qKxET/8
n1PG2PxvCkEeTzbA1T0ViV6sH3pc0tSPgTwI14nTOweW8U3bpOwZngpkSddkV0+pVjtkAfwCPq0e
6CGbB7AdOuh8vQtEQWPzlaPvH6iaAH7nY3bg5l4ZThZH54C3fs7HUvIOHw/8orV4UgA+oVlfV2sh
WbLO7t9VNwCmxcBbUdOxspe7R8c6e66IFbBitLpDv1JgWrAfBFdf6KAmzRMqU3pdiRb0LuU4kY9x
ijhjuF7hjC5HavBxgxMimeKrX7tV6gLUw6cFqAaaw9RrV/UxzmLllX3hJi7hcwDSIfKo0/EURdBe
2aicp2OlxgAU/mKTlxfAZEO2EOvF84YLyk2aNDPD2tt2cdIQwUykNWODPK6xQcHlKwjLib5EWX9u
ju6EndbKq87zBKjLIHrcIXGvbM3xZkmiOGXKxblsihURnHVw3PBhq+R6eRI7itZ9f5flNijRoZyT
YfhANi1DnmelF0H+C4VFbz/NOV+JoDj4XJjrTpiji+XtEGzxYZyw7w6DK4b6CXSdpMQc+vYyWUTY
09UAKcUqBXHaTcqsa7RKdIOGaJoIoaAHMAyvBgfKcOc1X0c6gtO8V/BantEI5pbtw+frVPrqPTqp
6sOWUoksy1AwdcymeZhANwzlkWBkD2a0bfZjtNWh+iE52qHpO3CusOWiXcyw8e+AKteffcc5fIzn
2wgs66eal8wP2JkStBFA9ySZ4mx2/SAPifIkDqriSvE1kRuTmTc7arWQ2S9oLy8hQii4Rjci1Cqo
UhZ/PX4fA5qrdjFx4C/6IQ7uaiquarkj2fm+GeHpyi18Swt6ucT1EgoLlaXXlVScT8RVWmIGUkMc
8IOVHv/FComrLmWANAUytYKv0gLS7RWKHe10U0ChCHC0O1F5EgjfSHol8AHDPTLHLkefwSUKoxna
ypNJAUHUiFjjrSUAykJjCM8jKS68rMs+YuNXeRx6LfQYwvLTc6MLpUf6lt8zaRZwzrHzGFXkMRoD
mYy/LSznNf+VMCRRinfDDrLpB0dY/bZ+t2Qov6naXE1qC22CCUKiFpvybPqx2bXn/6Ld34KBYlyw
bwdcXYhpXNmOn89vL4DPJ1RBE8vuhRGDaIhrgS4Uei5qDh+bdxl1S+iPluS/m/+lzDKyh0sfRCTO
GwLCHILbR+ntG8mKgTzgjo9FLNFTZ7bFV1fqHQ3tcuvQt5KEdYYAQhk16R2DmanKFHV79+WmwCWs
I4ZOgeS1B+4HY4ozav4NeqZack4x1hAFB8ZTThV+LKNXRugN/pvQj2SbiPwjwk+514C4sKUNgmaG
NVmUY5o/q/VPxqTJOzawOUVrOYpbtFYXbk/WM0HXzabAEC5AgXvQnPW8kxqvIL7fWs3MLZpE5ddf
cHTvyGjU5qivqW/3I8t++XVUyIpZX8k9/xR8NtkVd6aRD/s3jefzr7NWHKBUwfe0baqutn/rb0jb
qjmydbi6H4eM+HnH38BkRB0b2eHVdDjWssxrmLMtKb1YgctoHuouxJFMmY8A+GkBUCI2RqMGqE20
wtxZcQR5zQuk04OOJ7prIG/ZRLTbjKw6T0nVaemDj8GCebYfYhfOvHlei9NnK6tyMs2TdGFMr/pH
1OYhUV/DUC9DrEPfBAL8HZgwGWtrbaapZ2dplmysVD1LqOIOZJwiID6rHcAQRtBcy/+I27zHUfST
pghYFLhUQkm7ECU1+4PZdVmMnvWeuiZd/mhn2oArHDxuGb/Zr2V/LMiAIC9dl5wtiT59Xz0gWUsj
/UCKQVdr2blMlQgMvSwapTKZAt+sSDIP3VIHcqmjYJ/LjtrCnw1je07FL/zuWPungwhqyLxfnSWC
IWKF8Ft6u+UPKa7n8ZxyTGjJKZqhPxQXCpMB6+1KzjUYYudcGxpTPALNIwQ++owRJpGxYGMMy+7H
4+PtG3ZzOLvjobEQ4UtJt6nZy/KAZwHWMQNKUKMLe5X014Gh8ENrgRyN4XKlxi/fcykVYHChf187
4JdbFsUfpRc7S+IBUr6zvZOjuaxbguLFhkncocHl2K9ORoXNGRXMBQQBrtfPhqUsaOL+SXRYjz9A
57izkcE9oPL2Y3wyWcU2qMSPx9x9V222qgrDqVpOPF1epXrcYHlFT6UIpuXn/glSSDMVpCIsz8lZ
Yb5o04FvLwqI4JqdWAfy6pQkbloyuwYxObgMJys0Ks83UGVLtAlPF7qCTsUpKe+MdbemV7aS8UOt
yxLN2IqwNcT3C8u1Q6fPFlEw7vwyFsGrQqEZCnjZgz1aX6J2QBlSpMb9fw305u2OICjlq1v1QxHm
F8aMuJYq3jJgW3RsycoDVUxxvvbkBhKcy+u29c0Ht6oB9wFOiPTS9fLbP0MULU1Xe5P4TbuZVkeV
l2G6IPjTE0Vl0eU4lqbv4a6Dx2ZeHOckefimkv+pkoPRXkH/6kE9X97JVF6TDLW+NDMOuAQ1dXEz
SMdoAz0Ag7WHPjLu8aq/aFLccch/oa9dlLo85ub/P3VrD2ro0ucrcshQ93JhnXvXYHo/+AfX3+4p
btqTMt58ei9GOj39M/eOJVftNOwADsbOjQofhiWPzk7dvEpRf7JOv8rnp7cVAv3eFDEg1jzbjvSM
jX/l8iLqeZnDnRwqxRxi2QjttnTQtf8ylIN04sjUAVdJkz19pLFcM8CzMYD2LE3uPEAsO8An9UsR
MO6dXVgM9UEqjgP9QG7SM0+w0aVv0VFICCqx0NCmQfZk25obGOnTacIrzZCHr09F5NauoUpuFwdt
1284opyjitvaYnnBZz7SlnZvafP/S3lnYlj1j+YdnHF5vxDfsR5bPwdwjIxjQE1HnXaSx0EDaYrC
+3ET8DBkNq5RiNPFDXOLpAlHQoU8HptMvpib3Y2Oy7xkfTXs59GWyKvBFWLg6t3XEgfAFvoPUKKQ
VjR3ryFqWCK3GLowTTibzQPua2gM2N123DTBMpgknryxm3iSQsEfinDNaUtR4oZ6pNdClRGhUZfY
6seAAxATyU+497vbsNECvNPqKzGi3vIatN7N7vNwxStaMYDcrTvYItPeAQoRismjMJC4HWarl/5B
cPxpJDNcwbvhul9vQxJ7JugLi+yDL1wH7mX+eTe9mvmq7oEr99RRB11yQ1qQ9abyOY59KpbPnxMa
FWSd4/39V38JdY7l0pEUvRQ/LDpAeMU3sWNzxbE6am/sCtXdSHrKdeEdJiMahQ/iUqthraS/rHrD
P+PrRmoErOLePbjZZgdSH+ZxABn67/Jt/RxANw4rwdCgdNgIaVwFWt8Frz8e6sGyMw+Pwj16A1tE
Ei6jgvgYqMHkGg/UOzJzVlq+K3HsC5kaxSUv3fEPDGW8O0iAJq08ACB1/mQG0Ol7IOHxGfTBCTOz
zqZA23HnQcQeeY++eSaHjUZvsDQtD81OaHIWzHzNIVbUwhOaVcxTKE2MbswCIX3vDTSyTSoAG88z
zYiq2Oc8s8ffq5EFrmT8+OJiQX6p+NmCjnkh4iAO4WKLojBzSvxxNiuf3/gMTzLSLQ+g+iN/b8Pd
siAbCcvHRn3L5qe48VTGXLqXAQTTosj8i2iomlcMoo5kfGHY6qkxyc1eJfE1MTtDLNs2as3jhGWY
YerTjmenl4gWBNEmTjEZYHuhiW0wSDkQ+FxTt7N7sTSWh4uM4kCMv0Gp7R+o4r1BxTW07dIliEL8
yt8a9SjBANbP094MjnYUaMFtoYi2KT9xK9dB6jRDcjXLpGdqpxdw7f+KHh+3slNuzPdBcz4znflp
H0L2s5gg2/W5JIIniPgHXvVrDQgpQ+8wIm7SlMCSCsUHUtH0MC3gcBTc4Cp02ZoyWC5hkeZp3f+A
CFqYdv8GU2iVsF7JzQaqBTkAg0YeW6IJDsshLfV/cFjj64KoCnnrqf3HTbFt/FZAXHeMrbbHApvh
Qq/p9kwdDHndZ6a9EbajpB+QiyTfP460q/xzq/KGvVdf0CMf1k1AD+xxnMRky+CA5xDcWUBXS43W
hkRh35KCjFEm6YfcW0R87vmGSZGGUFNULg1r1mKW0+2dyuSfBTiRcOVg41gUpk5Oc1N1eaVVo+je
uQ3w76rK0PeHxztFdkn0JEGqodCnjGwoEeGDvX0aXFRw6J6chewBiUFFjpK9NVHCL2j6r5/lPv+C
C7m/nJKmwL32W121U9SKL3zWee3pV6/5FS2YP4JWudKYnB8PNHdEhi+IJ/p4QDR23GrvmifOuq/L
cx88B2MvnvgMjKCllUSz3I9i72B+t2S55Edj2LmBOZKYGXNE9ALpphQjmL5ZrAm/FZ574k3CH6x9
whnaY+Er6nwuwJ9pwX1x+jr9J1oZ+gUBwRkotlGLSsKyThNr5PgAPHQ7cTrBJYA3egmRG+juaqms
B33d4WXVyfAF7hDYlqSF0xIpuuHsg+2GZJeaWNS/7FjfnqDcBv293P3JjnyZLV2UzEb4whzMV9OB
twfYSbUnt+33CBqeGQ5js/rrdVTuTs3gLa6A+ZE/U2o6pqNVX68iMr5SR7+Ga55scHinKYqpHtpu
cMyfO/o7Gz03vK+eXcFo93HjKv+DsSLapLYywhO3oUrN8/rlRCOtFBvrn8f1G3FkHUt0NQW83+fK
eCZGYexBGRhgTeZHGIrexecX6A9l70l8Hr2uhPeo5SBzT8lJnqTy5OKS/2R/gRHKPDF9AfuR+5Bq
FeWGM5eEwG5VlAhF7tPpEiysZ/q2tRlk0zMurE6Wc9hZ3iDrA33ku/CP9roX1KfD0/MJrDeguuOP
+1F3FXWX1GHycMEaU8PLwWA2h7UJXsmYPHEE8fI4BCtA/yJzDseiYOhs6DIvCoU/q/DgyWfWKbnE
mkrRwKfT8s0wcVzRDj8pLx4b4fBr85VBwO4cnBDoVBp4e7wxOwugVMq3eWTryhs1o91X9REFjD2h
POm3LumN6SkS280t2tB1+dq511npdMf4vZQdS/60fnNEvz/tDq3gKuKt/wxFYi8emYjgTSiGlxQe
kHZ4Y2wUdYm9zde17Flzu5YMGAAxRGc/+324kftbrs2p1eTvkRBiIfW+F7fyhlUqy9pxO75JXGzs
77AhBbn+2QZU3XBQxUgjK+0SR8s7ZGlfPbqftwfW6ZuSiHHv3IIdGCGtpmC3MdkyTDGX6ICVEEi4
ShoeRQ/jgn9d2tM67RljKZ491sS72TlrSHJZILSVIzpdeZrpLgWpOePw6jvK2LwdrSi9/XcIH3c7
nlWDM5I4TpUWXa8NU7OCKxKThVV3HyigQ7arq6L1eQTC/r8w+/RUH4vQpEAhie+eiRBBDBsumW/p
yMpvWqWe9VNXwm9uw5ORIqFZOV0GWmfd021VRlpSlMVM0J+4l2nARtcb6OTWf+geabjBr7qTEbWf
ka2KC6z1fa+BlqEKgrunAALKF0U60PjNDTeTDBFwjiCLo7GDQzvC30WxRf8yBHl6bAOS8QGLFl1f
iLkSB9ALQY29KcNZOyjpW5aFee3mWLKpPIWNXj9YlWfwTzElZsW1k4oQ/XGjayP2mhZlxmm9JzX0
TU9sQb9+6tHQvxjD04IE037gze0mzzduSR2XgHhYrH65T0tNZ432LfeNEhD11/2tS4ULCHLs+XGd
sjd/FdH7JOt4RnPpGiQDcn2OVFnZ+ZDJ0SposoktHXJGe4Sq0GKNBKkb26BwXtrcxRyNmVBxsvVz
Umce8mN3eItkff8ZRH/2MnYDXiKbNH1AovA2y4NpI6lF4cB8dQKr7bYlg3fdYZfKKe4IKx5LYvli
VnDLq8ekigxP8cU/5QUNZW2oHcgO4lWU7ZWBjvGUzleV633EHPtB7pJTSqRIVOinAsOuz0Qfet2j
XLdtbXZhtAJbnAJy5Z08hI6zDbsm7e5SCh2E9vVyGglqppZ2RtTauvJAdiUtmGipY3BeMWbx7Cvz
iy+dBssjAgqgJjQ2zhPRmzGKm7ui0PrjQMR6dTz71pYPAxq6iCe3tV0PDLqWshYJXXapZmAXgkGg
7UlJCyjKAqp8U5kIi4JmjqlhsBsUr65fZOIu95u+zcW1nppB+v7K6dTWSgOSPXiC4VamNU3cFqCC
1+LAGHTMTOGLfbVVs3uXmJ0HO7MPgwKTTeq/67XyU81Qwll2aMtrjCc7G4/Hpd6efVmkU++qUBFR
v3EmMHYEajVofB266m3mD2c5h5WSiI/4y2ccb5hpkV9CokFfzxHKJLXiREz55rAM7cKwnble38pt
qsGbSiR7F9CpjitZhcc0vLCsFMD61NN+YyQs2EATRxRWo1nG7aTDzaFB2Fzh2xBslfmJTo9ZYPoG
qXeiEiI2CpGYPQwEZcmG74KK0nlIaFOPHciWaNJHRtjlgAPGpWcsgyYxmO5YhrwKUOqhp0NQbdMe
5c8rDrppUua0XEKJlzGgm6QdOucXNSTwNSJzwBhSc0aNicIp1UJGAbdQsmjbffje2gillddu8Jq1
FPqkPrUwTktBxhHn95ftTIc5Q/AMxOllId5wmT3etyWz+ycaglhRHgqPAamyt1mHLRK/J+8UK+FC
mxBWXxumIAcFMSbkyu+ocJ3ZXDEMgT5OGDdtDfb22Uk50UFV2JVnAyVOG71uaMIYV7PCXNiEgrFC
ifkjvLn2xuyHEhTEkdwTjWoeY+RFoiJ9t4clvbQUbQQ8RzoJtMyHbYyqw5XmzkkHZmHgaQVimjOr
y6DKfbiR8wNWza8iw5tGzcH9LLzQ3LXDVuIHQf7NnWTs6MjVLbuE6Q7MSAglfhyMqid4nL5rTZEr
caQq3BVH75I6Mva1BYS/S96BqhedWXVHjCVg1fnTe4VbViY8PrXeB4BieX2/F66jROYWEo1jI/a0
RAEj13a+BgjrKuVYGf4bXePl/krmaWIKpRd6OuWl1hCLyymYMF+9aDHaMpDHzp++PbXP2G0+Sard
bJwpUQ3l5FqMTGU4Uj0E/7yWVZcbpaNHde57uw9x+Y5fqz+f+vyITt/q1Nq0spE2PohkCq5eZf7B
pSCElEHRUbUyFB2rKXga0BSoX8URN4vnxt5gSaWgDITaJuys/NxwTzb7lwG9Qg5I/db1kT+D33XF
pmnsVjhtgTeDoyN5WjgxZ+aqqeh1H8zQhA2prtBugai2X6HGjjOPPmmauQdM+0m/cGOCqTIXdO39
jxjnWN+bV5v8HMzWl6+jcjFhK7rBcDBIQDDvQjFadxhNNjuThrVpkl6ssOXs5UESEmF/hhICi8Kp
CwE4u7bQUH0+bUMzX/XjpOxuIT5kVOHVCDNfKw8jrG7SWbNciqaOIpxkrvwN4CJv7kHU8WZEwSFK
S6r23DmLGh/FpN6LF7iGeb0tf4FUmyVXCX5NyMOYIYUAFUp7tCeonhMDMU571Ao41PsACjHq7i/M
HkOUD1qI3j4L5JxQ+GTAgw07R67n3XmOJUdv5eTDnPtpHBZOY5+cPpJX4y17Yeo3r/LTU5HUWv7k
EJQlWT9IsXG6s8hLqIrgf4rOZNVZhkysqMHacAxMpwhM6IoTJcV/hnfFMdQvKQFpRDbqRfIhl4To
uqLLcgkKrURv9bo6cwyYGPOhODAK1jrkN9iFsfIC3P+asuCuWcboc93/0trQBxoDcLs9ooO5NnPi
NXYpcxVk9E35FpS+3gnlu6smtbGMxLfPYOctymmvmtHWjGZYJZwKX2OwDAfaZe9u5JMK5xT1a2TE
aywKLjJk9QAPL4AplVA3EJpH8b3FHrtFOvxkMUDeGGkwOEFrJk8rz3ga0FpTiAfioUPf31bZvA6+
fwOa25hvyA/Gi6nKCY74AlH/E2+dzY39rZCD9dszbd+jJjBTmkOKvpLkvVDUuGx5bjSsNtkAVXqw
JUJV1jvWuAw+nnJfSGv/ViN79BNgGc1U6MQm/XsATunFayXUh4R+kTaJb44jlKlB7zJlwBv/zgrW
ieFWkw5sXz81FGdjZjMiNYfK5smSt5M/rVyCJV59l+WVw9kSP49+GijLGiE8pDdH+y6EslbsmPx7
c730eQlbN5DY1RaxOQQYiRLgxC9/0LCB1lMvs6GbaCSzpWrb//u/HuIhVvJjBL52Zs4KA/JNGjAf
eQuH+WPkRLufW48x0Pu7QgUk1uJf1Nl7KzELFY/EYY4ZhNNFVzsxJzLm6KKTu5YO/yHNXJH7qzqA
QS47ozBdwRRgVqlYkqGUHGlorUVktFcIwC1NPT/9SrPwCFbeiiLG9NJMmYFBehbP/JQhgU7RHzbu
LOiQa+8yRnZMgO1jmSLp8H9oy2XNi5aQpQacWmqiv3Y6/K8gxEkolWcKOp9eKkrOIOLN7qhIpZ6f
F9tx/eajfpg/Tm9uVyupXU/eLQ/Qvq9BvAhy43SETMq+ewt4SusTTHbiJwmjffs6R13w/ZF4ShhX
UvLDxGyjGH0HqCe7pxV9FLs3M14XE0C59aAUEkMt7WlUcNS6wJYV/LgbWKVkWHSZfXEN9H1XyYTI
b8JddS1x733YF8M0H5lckaguAiHuWMrL+/fylezG4yZMm7GZppMb3S5HeeB9eeDF/gVA7uOEHHYy
I5hUcuX3GKk4qtby9mudQ4RILpBcdZwjKo1g1C4Zk1enDFdeaJvSoPWFjx1mSWC9z+wLb/zeHuYR
rHWWfTwUFwPW/oA8qTlRJlP2nxMowobY/n+vhWz6lnd3G6hWM0q8v4ptLcONzmbDLVyfChIr04Tu
uKl33NEChBopMolhsLnUe4GpsCZNYDA0XC1fy6wMvwUl07i9XTYTYXkhe/I7WYi+JKE87EaqVbmz
g4+PQZi85bGo/Ie8oa0/1R/6/jJppIlt6JnXdTSPQMgcPiPbLeeTVTvv9PISia9tcAUaWYXdXY65
EhZVZXwA/5eNY9RxHBxlfED3bSpJaRdnJDXR6C5f9f1sjdmOyiQwyzJJyqJ5JQE1g3TR7F7bBh+Z
wEiT9JW/ectXzV7sPtPrq3I6kROrnU3W0nhN3orNrQ82Lv4/U1QHmwxGRDvWeJoSRTOjkGcPoJ5V
rDv+O8tRKRs6aEQEPKGDsNQHAR7iC79NHhEvRgQ8ykNiySe8EsIyBcoFtkvHQq7iI1GRFgVvVTYY
RJk5jKWl7bg+OQ75I7yIIh4GR2EUm4zrzwRXt6VrK3gWbWB5rSoY6trMy039R2W1W0ICLPDqvSVL
a56IeMTrtJHb5Te1Ko6UWeMCEL5syFP+5217BrTnnVGm6blROkI6mltNwzD52BG4n6S2bHmJn1Ng
0u0CI5W1nVRgTK1WOBF71tJzFzGgJ4ptfOkS5OfFADMK5Q9Nluz0E+qvVbB1ASXOzvGZY219/7ib
QgYKAetiaqSZf8iTi0vzNx5XCWq65Na0sjauAawLbOTUjqG/9cBw8G0pZHjOOkybYDQrHK/gO2lk
r7c7c6ncHu3gvcgGz09BkF7Af/0qdyy1v0XhBj7FVf2aFNGtJObfrZkOQkq2W7O46LYuT+CWc9g8
1SXFu3amMoPf7k7/FKHiO9CSCNAqq3+QVPODX184MdXrJP6regOF7yXqInMG3OzRzxl03sJq/vwM
MtMdGk68To9o8t5U9uM2dYznSgPbSSp5DQj0dzuUTg7YWs33saDuwGTq1iud488eb3aiF5442HJK
7U1hZnQGZudFyCZELc+Cpt2r5Sw+vy224FMQyBxARmi5hwoxbHhTLFgOEfQc0gqD0VtLu2TjztTN
sVi+mUDZJ6hwlWke+LY41Aclbe+/5q2+5l+Kn3f8Wcs3h/nujIs4TWgviFKit+/8Gq45JOFPF0rZ
cDrJGR3fx6hCEyuGo1dfBPEomj9C5vaUd1Y1J9lRM8+R8uM1bH2glPpmBthUN8xRhXOvHeKMOKVY
dYQipD40OCAy4mmhwbMKnSHFxL0EeG1rqFtWmLcuoiRIggvfD0sp6auqGzqlmX6koAmzaQbRthUe
w01iseH3zJPYBSNLOJxp+OkStPU4IIiF185Wa8O48ouVHeeBWxqh/0ZxW+EMa/jCEt+WDdImLw8Q
du+ZmUovJkR02cK3/fYcDaP6SdvNV31tAov3KThjhwasRazmFAp6wpNU2bmsVsf82znFivYVk98c
p57lxHDsJtz2zOhdtfvMY1+FBdKV4gVcTOeky12dN0J+HIKHe5VI7fIQORuBDss07KUjRhFWCWcO
JSv7SS7/g/2MKnhZ2mNSAx1o32ymaFzjTmd9crYvYYnmWS1VMDlLxV7zC3iZQ0s4q1VO27rNBBI4
CJOO+QLP0792A1PsAcLr5g7V+hA8dw6oK0jRZjmifPFugEoVbjgMQA5j8HU/9Lvd+Ihw/6q/10s/
46Anhu+mvBJ6/YtDMe3ecSiseWmGcBTtDoAl9LlJiIg+JenyEihzUmDS+g8wVrTkBT5/ejeb/MSf
NdsuytnltthDu/HqyevXhSS1f7Fu+Ak474fI4FbdyYPET0ts8+F8OjUTEG2duM2bSKSuGjTqI3kH
aab07K2/WNntdWmnGNrbNKVFWlC//n0QP4ACqBa4kqjrvVsMo1ngS8gx2zHoVJoRy95T9VfuogaQ
Lv0LLWSQJ5F6fJ7AYcTtFLSuMRNU+ei0u/tnVlbLzh2uZZ+5/vY6img5P3O7rJkU3+rgVWx9J0l8
GJbQlObh8WOvwlKFKVXllETBM6FIdHbc/g8gwX+TV1Mr+/MJefFQ+D7P7atbMLeeELV7mUMbZeX7
BAkDYhzFOfizJt0rbyYSwYkQ+/aYof43lRFk4K6re40glBckk7r9giQD0lY1uM5TPRIsc0eLG8Nj
8bzTHSaxLDqqO+nfkZS+r+sMO3H6V//vMpRmaDi8sII55dYkKRmnrQ85gJWHYueZAGe8jkIS3mj4
fDnOe2traurSLeuPT3RS2GFmkOZQhBxIddr6ImBolhi6iKUrTyUyGPv3cWnVjp8/QbCqcOydDjKk
Q/b/7z5A+OMiD7tNiq2v6K/0mEOOU6mNwIh78lw46nIkXoPep0CGL8UPA+r17XtfbpaSltVt2V2+
1CCdD/IJwR5WcMFPwJFrmA27LLI1mzgFCEwNSNwNt0HKknogZYlpIo+Mi1k3U5E+3nbhPTkauOBS
OT7Wbs1XF197xKCNetmuJdPLHzNOMvEJIrEtzkYSMoRqT9k6AFdUCdtYuLiFBSbmWpVmaeVoUdCP
CprtNQJAqyPO9SbGD45PLisjiWTa1hYjAA4xp4hOE07vJAY1z/Z5M7pdur03C7FrE9eSrkllnuB1
1BaFFNNWAN8pHFTg37h9sVh5fNHRfUNhqULyiMAQfwPdk3UeFfEr8hkcgw3K16XhEN4NXeWs5D/n
3CpB/q+wl5LY9R27sQeG1u3m5VOLBCBdRQZtblk1yrL0zbbOWirjP8k0jZyS6V9ofU4TNjmnaJwl
KSx8iO9g40IpGc0L4hDeR2dEbIIpyIzThZqT0GKrLn3cqWMtXOVk3BJFHvdGbkAEux1z3mLHvcL8
HC/qkv+dcrSybzIe2GTZPe3qqh6bT/YkfwIkLeTnKyR+M0nPHvf20Inb38YOiNQ9q4sazhSUZHMW
0AzM3iw04kCbrj8FPJ0UIyG/WDnaKtQDrEKUZuwCu2Y2ikdYgKjcnchI6EuYRPUQt/5kbM/CfEAG
yJ23HBS2vWeUH3RdTrh4yGQjGDrx0rLVyPsUpj05Ma4uMGjgMM6Wx982rWKcXIaVobXJFKKTxvcF
m3EU9ka/M3e4ApnzFwPftqnuaTSeluovqQAAA7wsfTGD8m5wxVPpjVPnsz0FXvJwg41QWkpWYzZv
/ilCg4FD/aqMeq5DsQvM6aGchvho9XaDhjnVV+nIM8zU5xLj+yy+r304ya8ttAKPh9fFnKlI6O75
NcC+WbHy0xKuzAbYLQ9paYtoZ92hlgOkkuWHINbHKQvKkJA0r+nCXynL/81f/+L+n9IsBVjynwI5
vmbsVabsrbwstTEObU2zEzCWTMrv33xmNgDEQ6WU2hrtMVWImyziPmw/9pwvbA15xeBR0/f+kNmi
Ra365i5/mumSbCBszrOjgFzy5wKWlQeQP4BtykXjh2Y16jmT621SOGYilQ65c+bof4K5Ol3Mwu/U
DxnBDj37ukDHA9vl9oSNtTTFyG0BM39XMW+aP1K827xi14c3dv/6Id4iXsTe3h5r4UrrBIZN9yYE
8D2zP93X6J99SWUcIycVDb0sVZJe1EIj77u/oWFxb5VVJAmwmLFeW1BMqQrGSmhHgxi8tIsafLf3
zU7vsc2sSxaJcw4V9LlB1TTvtYVD5X9pxvd8mYS6irKAtAd7AXhJHCcOWNPDUGz8asB5hxsABKM2
bL29bpzV+pVcK/F8GCDmvt0QW2SvWBuuDK9yQONHqIP4kWIERN/Q4NtFijNOPF3mTLx8SeADNhfB
Djhnlwr4xZ90DPImqUtS4uBotxSI992xLhhQ0Mynk+zwUQfv7FrcaElOeKw0zzYaybPi6vJ3FCnI
K0oYPpqhTo439tfgcW/ZEw9V2Tvfylj5vAOjUSAr0DJAyiNhqF4X7oWXZ3xz+xHNoCXBAbL2KmFf
L23E9EnFuwFVXRx8EcITB+qpthXG38LQde6zOgw967YPvd/pvW/6h8+v3GRUTSDeAosI6g2aCWML
8nDOHU4+3m0CcXv+wokOUWkJLdrBlMVKX2m+OUN7jjudkD7u6WW1/kJ3h+M0GfXk0Od+ew2h2LTr
mE3jbd81suoKuki01kHuCGf2SllCQoMqYoUVNcN8f/NgmB5rhpiJ3bW23qGzDoCD6zFrcMxCWRoD
dBP4fhx358bRldrmq1H0RPUqWsX+22tnJRuCuMyVDmG9k5Jhkz2f5R/R72q9+T6OKZ6hNfFg3pOy
3KFuoecicg/+GqSVQ+cubMFK3BtW9TuuuOLgQxDN44bvhs76TFgPZPZ+/92zpY6tUV5jTx5ufUoT
5N+8f43Zb1aD0LSVfqRhkFro1QgALmw52cS2c5Vnh6Sxb+aG3xy5UEqtXlFx0b1CJwvqKMMEC03L
hQTPid18U7vfPdpuQC0XhPjZ0pnVKN2X+boLg4/wFWaz2xYV/QI21edqORe2Pq3A6ZWQXp7804AH
gOJ5LDx3aBbUes/5JEcTCI/UTWHDuuclOQ5oVTkRXSP/81AuxnVKqU/yzgAvjwjvtotF4qr2F/LO
DxkRjqRcz7Upn1EZdjbDuvsshDf68vlIgdlm9eBKDiOWeT+QzzBN76yV8wI6QMdIsPzID++8clpf
NkiaIjDGF6sHDlm1jsgWsyBpYDpvErZkbHS443P6kgLiu7jCMil8ODthXCt3fILKLXn/YudWbuQL
JZSu97x98F5qKPIUkgvDxv0lsyATWdzKxxRrzCAeNgU3X4dPWCMu3Ds+8bpO+x7orKUd5QoD+yci
mZiOGEfKXnkKnsO8fcoj6cBL2LVKK+GbjLZmUqKuvkDAk2HdVjRltFHxY8b1gzkaOjTtFXRPN8qI
XrasosiwSZbuURr97zi21j7q6jLAghROhEv4uR9tRMUcQ0JJep+nGP9k+DgDcLIPKgIMwOQFEFkt
kSNCdXOnN34vzFllVMovmpAar0B5Mg9yOaNUlQAHNmmziyeR7zpa5PKoAsZkCGW6LNbrs7kogjsZ
ll9MHB6aMIFibBpVcoztT/VcPYsfbu7rTMD1LjCuFURUN8FIHxNhH6KR6KL9b7XE+5V5qJnOmZeF
sclPL6SxOT8F9iD/fvA/7gReYZD3YMJABpL+5PK6KUtp+Rfd5g4rWIhGjhY0WTYJhU8pprrn6hu1
k9nC0xczFb714pXAubOJsfbvrhDr5ehCziP0sVxqCNZ2+S9VUyHyfhsdw1r6ZrF7LlKJmpvNpNyn
/CaveEfk5SkpT07nGFInPxfEdw0bMAx6r2iIDlTJiIdNxCSNp+aJhV2WylmdQdDYkMLKvD6NAIQU
9MMm93zetZfTi+1ig81l4Go6wr9LxDPWTWj8W17WiAvSwixLwl682D/fGxf/72HjCEVA0HIFxM57
l27uNMIwj4l+DWNjEVjCVo5kt3KgHvoB6zUfM5FFz9zJwZu5xqWPCf3oUOwUB19WzqjAimEXWCor
3mQForlPw6QV0O/XL6RROy1W5OHVOEZsLjJ6bfSnivecUw9UCW0MH47AMZEkEQuu0+VWopGVzrER
7CK7QCwYhZ8TWz9FzHWMbWdgMLVAmsnl2ZkiUODJn3TCLcQzkCVEWcGL5aeVxcamxSN4Du8dT6t3
MaRWo8V/QtEuWYS9oDdQGajGlTtsUZCnGbjL96BGtMPYpwMvcqbzCascdGtORr8RMYo+DZT2fPcr
9QRO79e0m8tuTesThBrhtVz8mtYy0MnafU78Vgp5dXPJRyl6Hy1vM+VZekOYG/hlrMaMWdsBIMqG
Q5ELEzV2r+CCTdpB8uEUG5zC5QvHZKdVep9u/8dsVDzwYjQZnoOYpaDa7GVldxG+Hfgh586vPiIq
tR83achxHOeg2CRIiK6uP4MHvJfE1Mep0h2WEEC237G/3FJc0/Mt/m3dgWvFPd8so623FZBDcR3s
OhtIjq9BiMlfZcDc1+kTUHxjwI3aJoaNMhH3wD6++Mg6KCRMvBJBnvLB1Xsvc2cZSKLLvFV69saF
qcm0CLoXc2uPK7xAGDdFbGKwvSy+91ZAIRZX5AkvU0XkCPc1t5XV6t3JUFxcu5S/hVOaLf91yhbe
q5uyK8iWUFlEs/e2O+5Ooj3N3gkaTIA01M/Es9Euot7ttwP6pKvWE74vzBZ1BpJmY8n0IFeUOGSq
gH9RAcIFgbTtIjqoLTdifnAqhvvemiKL/yUH7eJeQQT+1vrc9CD+6ye2mZGuwgPDx7akvI8G3c6y
mIJy/NntxSyTOxcQ2ene5/IgQyk30660h6z31FTmaw3p46afBQ1xxYGB5GfqjFmK7FtvpqZAlUHJ
5HsLA4fPOzv0h9AQtVsRkmJ3SGK1XMhujF5A9xnysJXI3RQWNS9p7om84r6oVXtmAxOzAUMDH+CQ
cgCvfETBWcjJ45+g07zNaXPtLaLjbD9RyBjl1yRcBtKDglSG82zGm0/BeNDK5uo8b5DsXMg2vIuJ
8U3mAn6+kZRc4chEItTg3Tkffbdq5hRzLxPZbS8BfcR6uE3LOLe67I+nsYb75lagtxJ+yrxg2Hjb
jfHzpYV0dBiyQdnUvJoK+NSwxUbYmBKAkarWOTai1syfyqd0IzfVbSVH8n+vk5axRkfN8yeAFdt2
RaWyMs/UW8B7VvIVhVTQtXww4CG6hbb4Kf90uYL7e1r50Wxy3YwalxXTDVUlXdHm/LfCU1LQyKMD
GlVZhvsMl9amOlLAUi8/NajJY3Pmkvf1j1sVAzQCWz0w+Uc7tMPG5aSvzgRAtvKjkbs+FHUE8+Vb
NNRAVkiOf5rooCpYC+/HoJnxqeTtQZpyw873MIkyhBMIBv6BMKN46SOAvXeazI92J93Kav81Ywzd
gja7Ea454pyalk8/zUczsaq4XHscSd+y8LhDqEELemqfw7ixt0epJw2yFMBeoUvqeX4qVQ02C4qJ
Z0x3NfgWTOkBJ8kT1USw6iN0jEDziz+mIZVe0JhLp7+DAQOaUyr+LFsbyRIFiF0ZXw/NXWkqGlpj
RFIUmLPZZF8MkA2R1iqQ70UWHBxlHS6oLzztyISNzzeJ/Pz3hYlqZhoWXFQW4SrSc0ucXmiP/uSK
sVnLepBtrMfxryQ/VXE+0HKIfs5zkhuE4LsQtxnNmcPgrdBIrFAIou1/TdNKCvB/rknOItdXqGqi
NFdd7g4jV1rxtbVyflrxToKqOI6Ss8h4WYtgPhM+vWzTQWxxZZ32H7CStgsG18QEAsAAUfG/6CFJ
8p7V9jBHnhJm40cgbrTn0exVJXm1ymGszrHxSsd57NFSfYMQgQqvXASJN0gIzI2uzQiQ49l84Kud
NNQv9fYCgIj8ZzRV9AN9YGb5Dtv4WUFbWvLZ1EBXLzb32608zhdHt1Uh+SQoOQbrgXAk0Jt/dflI
1Lqug11EjrLJRWW14G+UhLp2bgHxHWIFkpeDXsdkPZiiIVj/16jZ+isxu9qvZBcV3hGuxCr7AjYi
nrh/KIp0nG/+/9wLqgb9393w9QHp28662u3nddqfIqykeL+XYztzaXbVz0GdJu186tt6hEkroxHs
b1WEKbQCzQM/hWwdRhI8ijiS6koXZqV8qA0hYw5cYRBpRD1dG3quFYT0ffE/cPftgmTxoaFLzcoM
NdNSGw2WuL9Ysc0gpVfhhPk8ecnaexyIHo0yyZ8134maakZkVX8AlUTak5CYkZE1EhvRcrWGsInL
/rDvKK8zgkJtwU5G0reRu7jciH2yYUAXiO3wKczA+3UplONOAkuEe+gt44aob/k0cipuWYdonYzx
14aZHVddTIpnCx1RRokYdnKZPam0dkHQWnWthr8/5K/+wNsVG4cYfsZvwrTE3g1wfeSTHk1BDeZ1
gy94+oL4vDGsprsk1jbkA3iulWfJUrhrahD3QVyzNs7bO1O8JSRUGspOGU+RDMP7S6MCo6+9ilQC
LAC5LtjsIUfZV6Rj0QszPAZJ+LE1ZeZzI8l1nEgBVDa/stENLuT9nKOZ9nnECUm7aLBOv4VRZYiY
vs+oXRkDVFcHWjpz7fcj4HXg+ZfBE/58PrzhoD5S0IaP/fylUUh3OsZyAZCg4u4yhudOHmekteik
Y0iDAAJfLzWWlmmZZbxGhuU+tNnluF8yW/7dqkRxWPyKg+UiccIvF4xyFPXYulFF0gs0SpvWIPM1
MHoWCAHsvL0WQVlnqVKPQTwWLiYHLmp8t/gPhhO4f3uMgFmEaP827hpYUBBVqvDyibOOrQNUXEeb
n+53AfVwjykDVd/tQ/OF2nB71EH5R0Ulmn/yPIeaXujS7LaDeyVAAzxiJShthYiZRwcWoh/Hbw0z
3cK89ZTlUTObEvAGSD/aFv+3uSHRaRdhPhoaTZMrHBjfR26S1KW+mrPq1s8hFTmnHfucTXDtZgqa
VJ0crqykQP3DJOUzKaqVzpS2dJxgZcQ+i0A9JioaMGxBfuACJfRYrAQNg5dmfuqxvLP45qLotGq9
06olo+BNNOR6QpiERKdCa5T3bDiZ0N1AtpbXMCeImm/XLKfqADafvMD7+P/mF29W2gr9OUUWp8ah
8U1w9PKZTRxPxR6zgGJPlIAX60aFn+hcPtcMznGBLVChH2QT8ynefmGrOMW0VXjVpY9h54MGp0Z/
4iqY8K6S9etTUEJD7jbfUUGnnYDeiQGp8BNXP01l/ZHP4gqtwhhQKcyW/84/AXZrGWiqlVKAm0+9
Z1CvhNayBrB+HEHWRTgc0qfhMIa26d5vQ2NzuFV2aVuZZuUiUIeSNvBh1ZyB6gH4OWLydIk91f5J
KOsPUmVbHv+T3N0z1gHUKmhoSX5oX1otB+ja8DYbcG9SGcgV6+g8fRPQGHKt3TsEn0BoygXZZFy9
ANwaVUA/Iv89P/Qvs0h1ibzWY4yE7abfrcVhO8W5uDzi+IDHRNoq/zqzbITMLgPwo2GxrBCDVG1U
vjllLByqvkVXh5tvTfEYCnNgJGx08Sg0NY8axVxwEsqIFrfHj6M8jy5mtdN9udjGHCkPYbuZsU/y
lChnEN1Kb7ZwT2g7+7htmLGXGrVbJ4Fia1ED8KGwfMo1QUqQtfcs4gQPqjHADfqukbCWWMQcaFQR
7f/AcUvFyBhf16Aal1z6MQdL7+8xiF+LuBiBJAmP2uFDg0Kb63VsnOiQHQ+4l2yjyE72rX4UEUAI
ttH7BBBu/7zfq8CFquB7PB9J9YvA9wYU7q0Y9ZJE4vdAp+EjZShIC1jkIKjSnQNzjNnlVcNydexp
WFrYt4bCWS5vXhVwZbCQ8gAcqMJlD4ev9mUdcm6CmW+fi72DG5xxlPGIg/UTTrN0Q44vqlCJmqIs
GXk4FPWNoktObDU2aEcrOedTpGpt6Bcq7iokL+U+PPN0wnrLsNZkhKHaqSJaOwTv6BipUeH7GhoV
tPqE+Am8gkOzWnHKMK9zNVuqEWkiV91gCcVsOA4De29iKIHuZA5PSo7ehK0Q2cigh6mYiDhu7jLQ
JqC9Kw5yoUPmH2ZwIaz1/Q9DptYb/yGZB22CKoHaqO5gM2inah0dgsH/fbNzHSMefiamWnMdiOmy
yvLEdbjP3GWHPDKHaOz45V7S2E/xYpAEgld8bLr5qRLWwe8162diS2HV6dWCWhmrDh09+7rbvjAX
joJ/YhQsz0RRLdDIOlBewjh/HqeR+YaLyRTv2wF1HhChnTaqxaLSQDAc9+FzaBoGq2YPX9glZdtz
j8MD62AbF5bN2XEhYMOit6XsIiUwW/Xl/R2++F9QqTAzHhRD4jdM0mCHIXbP8pL4I5pBHWM6wk7G
QL4g4W12lr2yoWp9LpQg4Ac5C/vDdJ/57ISePL0uU02I7LEdS9NxfuD3NEekIdv+cLg7u/ZzruTJ
ChS6vH4tK1hVNUK2aMAgAmY8o4qkZBVdplRvkj0CGHpXU3ltlTu4THFXSi/nwDbaEBspMsRqOdra
4y0DO/w7nUGEVrzn8c5rIZ8UkBySW+sO/1CRGkEL7tUm3WNjvSRbRvHzuX6yNnmPJ6Dq6E0XkuUL
gD6gHQJt0xaYlfwLOon9xc4MSCoG6JoNmY72elF4Z6LCjbGulgMHMZhg416XfikUI6eQ+gbJKDqJ
cG4R76X3L8b4DwSOpBfVDOHTMpYUXneBapIX8+xAGb0Q4wj0FcT5uI3IEGLGABMgglfRUzzevSKb
u1uVZ1ZtMNah/Yo3v/l5h3yhyEmRTTxBE5jwFKx0Z8sTjWn5Xye7yCMhhBNMUJa0VGTd+9o0UMjp
IS0vno/wFqU96LBfUvCA2bB8QByldV/kZSgvQTEtvi37bf3nCKDiioNu9t5Faez6yg8/OeHMa+qs
i4nwg1CQYQZ5ZLxE54Vwojx9mvaRSquc6EX5/0MMk0fJDTtCFMghscPuOvQUPkiw9/S5rckN5Gzg
hcTIIDJjEcKhVBc+cFP+H0p7QD51iZbogIzlXFgA3IvErDHAAEZuZ/jV/prl1LpipZ2VIj/9NOlL
yKKrZxppqqIW08AoYKNI0MGIdwBAsthtUqNCB2Ufl+NmYSk2D0PTvUbu8TdB6o2jxNGgtF1gPdw2
mzbzg6WUKOVuD00sMhCZJgi0qv4GGSoRjcuxzM9qnGmN45p5LdZ1jvxTxRgNOQGfYleOj5ydQlbF
rL/C3Jqu+DKiMmpWEhPSQq3mEj7hgFvwZB8heeJ7R2y99mJD5pZ1nsnMIuqlMK84NwU5Ed5E94jK
qW2hiKEae4KOdeufb9i0R+Aehg5e2ogKnAONUoxdskzgNlag05jUKTqJMXIdo2mGwZsKGkJVlvnF
HZV3w1tj/ctomu1n3llpbN9Uc+wDz9Gqe3W4T/G3fHsIMJ1i4kSM6XrZU/eEYBKe2j1GcVX8b5+f
++aX6i3rx4cq1MykdOd02S7gn/fTp9rWo+eLVEgFUK9QoWSvgbtj1rHpquSOzV78wo9n32MibH0h
9j27uxUxVJNtXVoERjQc6dL5GVyuu8O4dbfKg0xXcwU6beGWss/Ul9gLnSsPyrFQUiLpdrFXYnvt
URfH1KyAIqV06mjVPK76JF3hchpyuobSdlS3N31MGyzKFwW01ZOwmDVygmeLiOt7NpIm1rChQ6iP
FHYQHZwRunGRStqFdj9acgKp3ze1HywhecV5xefhOvKcoAT8ewwPtmXI04AXh0w1lp4nX9Dlvsmr
YawAiN5bVTeIMxUS8oabcVA4nO0hNUgMlrrlh8Qp17IUaAXdgWUVBbxTt0/m92K0nx5b6funOkBV
9tLZGMxjkMSGR0CyE+o/4rbqIQRBPJoWrmiR4VlLn8iMaSmwcGXtKDHmpbI5Fn3NfRUimN4ZFA0w
sLUHq9BmJS+j79MaYYdZDwUem8LpCqSzySA3EJlSh6BAjAk4RCLGb6iLFLe/vZrndAmF6GdpBNmE
79VyMzvBoZhx7oV6cU4cHzNBEcGzuCu0t1akzpjXpErs18gpbC6NRsqeuaubv9AkmbeC7Z9Oosx2
JfsQ97NY/0mDedl9/CfTnJ06LfmhyVpXOlGYrbBLouUW5ZwBVyu12aVCSj17yQ4trHheutI2zNjE
3yrcXAvmlXk4JVDMuKyAQgQFeOYSds5/eVFzgWNtogQ37QZDK4cbAnSq/0gAd2YDpltI+S35kYAQ
KMvy2+jJDIOczkugq6gCVBCXgoNgD7hI5OOhgUo+8qO6x8Xo+HufBTusQY2wJlY7kiUfSxDOQMQu
2eJj/43Rbi07NKw+Wrg/monYp5ARxzSm3Wn1rFRZnPgDW3XSvugvY9mNvMGwwZ84LDfuSPaHvffv
2YRou5zXRT7UlYyB89d1XjKFy0Xq5nhzr1E0J+Irq9cE3zqM57q8vfqnZx/PPw38kP+7mtuEjX0W
re3fBdKGPo8OFeXD9B5kJlrFebyDe60VS5tGuJFAw2uZUdqWrWRZM/oFGtvDDTBRqubdvDLyuoYK
tn78eFABzWkygWXl+19i+qaaRZoY38zYSYUJiFaPn2u+UMgb6zCzvFs/tnQwJtnRPN9J8Pa9B2XA
QhY7UNqkaGgGJNNpmzqziAKfck2xJFJAolJc5XlIEMbk8IWFQXk8AH2do9qkj7F4qLMUIg8KiVCD
+BhzBrfWUAHp6L02FHVEJiAmekDLzJP4D1yA0aPIrD7MbMPi/b0iTR5bI3/00402hzf0P3ze0Vbj
+ruOU3IgCBZEMXBC8VIavM2Dv+mUOnTxxyjTx2vOW7aa+jBqLsZY6u8dzreSkYGNKT0PcKT8Wjoi
9gTl0vlGbYDQZzOonIvpJsjyNzzH3SsWl6WeMFDn3BPiZeguyTPJOiQ6qoXi7qStMDz2DTCn8bOw
7JMi3VJzrl3V3rynAYiKCqelLq6G70UAGAD0J1k5iqkjeDS1zGU6EjblrjryTV7QENRcV79bglQ8
gq/RIHu9K2j6KZ3mr9nCV3e4dWriP83z/n7nNtSgKlAj5HV3q1wdmyI2p7g/Wh2151SBCVWz7+g/
td6YoU7ilbagMs/+9wTfvgnYbKp+ZUwHIiq8/s3twhqRUlpq5B1szsOpb1R6hgjTFGfu6vjoYgca
FQ5reYKXsLwLqD19NWbbiYfEK5OccL+3x7wEKV/hKam+R/1yWg99wY8oGAlIK4XDkQAhhPP23pAC
bHrI4yKKOYDS5g5d2+bfnT9PadcAmFxa3es21O76Rt8LQPfwBNIDB5IqsgWneoWJevxQqmwG5Snf
bw2O25/rANHtheT4KrYRbbZlpASrsYv9fWKMjKO/fsq3m1kCaRHDA4bJu6HutWvt7V4JGeOcgd6f
fHW8OoeAdsypVkzs1Jm8nYb4oPhZKzHQcQJlZySFTjdsCV3HxN8K8XT85npbgRZZhqh+BAcB5L/r
5eGcJP61lSPYvR5UJg5arZ1yCoOpjcpB00VqDq4YqcLP5fpPlD8W8doZY0oQSw9gdgIlusDVL1La
B6JMkiPRZ7yk2aFQNLWdLqg5y8wzd58EHt3++GUznuE4s/f/DqeohP3tKHl67lHIjpjGIP+5dY0K
TXwL/d/WoM0FqAVwmojFnj1xVVlIfIZ8oSOygHPzLJAYxUsKmMZlF3p0U7qYu3k9XMNxrZ9itO+D
2yT37DL/ZSLWkyyEqojUTr50lPPU28Gl1dhlvxpBEbzqH0MkmAgq47AklsGgGwOrS9CMgTRtancC
WV7fBkPth013+ND4nD9WLLg+PIIwKDZGCO9oZLsFD9bzzomJcgV7BBUN9udIzzWQC6vbRI/98bKs
Ct8Qqh3wytRt1vQqgTzj7K5/Uz+/T0IKFfCBnElHbCRcUcAu5saj2VNg0LONVHXOTliYziygaLrY
7V4LJoSd8PKKBsjd1o8t5qIt75QLk/JVbxryU2kURR8+0xXdsVNUZcdEprFmD6UJgwWOzxytgHIJ
cLu+y0JZEpkQBCSJypwsCxeS+8Fwz0Wlg26ARn2a39Luq40uhtPBytNgSoms4c9ckzJyP2OeqOHB
yDKgfOSZhFn+h+V7E6nZsMtgJ0jfGfWJ/us/tFeJ0QXqPQra5yFaZ8k3jJE/wgZyntjWEgkiohpW
ct4KDUB6WkRdoJGW/Qg+IG1L9UCBhNgQxDlTaezBBIm2+J1749S4OKdhkjTpl4f7MBMYGOgmDaNo
YCwZDx5/7XwwTVLKGY9CkKdqGjeeXf9gzDgZd81JamcIIfxsgBSOTYqty/CUsi6aQyU+4XUL0wi1
jZidl6JeSeywTmgV3M5ZBPcf7DVjfrDEudZeNdN+/deKwVMCx6ksHcK/7ZoHt0bjbv0KoRovflwY
ADHyvAj2AfWDJzviWIExzAZCplA8IvzPdLEoM7RvLzTRnmtsTtaHmgrLyIuzEQmxddNXMT/hfGb6
Q7FDfpyPUOTapRu17fGO3braJkrG5yf7348Eu7QuFV+ztzyPnfgmmlZnbflMeKupub9iMj+92xKU
99knJAtiMLZeYreXniQ1MHmJBMDsjE1b6T/3dAr14axvNfVDOiAfqgFswQBWFEM5hP035ZBixkJq
yWoUVqFA0cj11LkHSsNd3XKo/071kDO88EItJzA7LKu2TK5Mpb0js4M7n9kBKw2Mh32cxeSxpWXT
CokeUR88+u96zubK/fVzn7LTJKe5MjMjewQ38PjVaLELaPmk7E5k6JzveMnv6ha1gqBnxdxPo69k
OZ7Ogj/z4F+dfdbZ22hGWnNp0I8sRnlxiHwx6np2N91UtNezWuk3Tyw59rI8uJNuf7K8DxPtpqyf
LVBjIl4aUNueZ+i5AIYJxI9HBWMQhHRVqmfHoSwmtTi1sEDeO2kSz95+TgZ6ZrdSgSFu7xkJWVS3
BAoKVSQhRAGYtqMaIXOuPe44uXXoxiGNPnZ8Hx2yMTMiap6tH99VYW2OXkPtqp422nr9aUuvCUqg
e9+KBGlK2QXYJaGAw1LXZ2Xztvl4wMgW56+3az4HObo4GYbc1pWNUeGDQiGhb7XEPmxqD/2S7x7A
5qR4xCJ1YNZrySkyCT08eg/XAJmTor6Pkd1ePh5zqslwYem8OF2gxpbkD8xDsj1sA1U1L1l+KUd4
Mxf5sO16xFlb3AUZShmmeN0V8dxB8FvA56QkTuy58/vT7S2GEPUE9CASFG+mtvNd/LrqRVaET3qA
L+5Vt6upw681TGlRpj5YWzicYQOJ7pQNaFxTHwZY6dCU0//671bpIGSnlcxh3HNeMiniznULj80U
MBlCB4qVFj18iTXbwp87Ue4QOTh+0O78y31MDi2NVB8iOxX1mB38Ki9ZMCzwvPeoshbE/ci7uix/
pd7a3IolSlxszc9+XtGCIFwiYr1PByTeHULUWEkiij8idxlZFXyBktisLgYNtxp6/FXBhiXk9rx2
D+8GYlZVjUr73k7oewzGNU8ADuxEPsYyPsKwLx1eoaNItp78envXo6PDZcq4xpLUiQLmn/1HPZjB
zuygEf0efGguCPVQ7bYayL0RKTj41NzrHAPHl6aI5FF4HCcumUoVDu9jh3jUNoSbmLPmnpl58+eZ
oe2QtN+py9y8dN+WBc4eZtPYii4dMi7cm3g4jJakU1Rj5pvId/Mk2Vx+JDQyMc0FD8VDyGOVmDdJ
8X4CCs3DV4zOIAKL2vdrvjX7OkLTktH61BvJfIk/lYwJE92XRS49ksDf55boH3wIe1Th2IH3FUuT
pMpTz8qoE5Dlqw+i2JrSuhNiVKg9kOQgnn3tWngSyweSXgULxF053mEiCiHI1XJxJqa5Qd0jaF3E
T3THpJHSjJbvuwafHRsk3Q3vzBa4wv4pQU2ZosfJyhamvytHIarO/v+wbvFKAu1YN+fzt8YGflm/
jBHwY9PTh5arTGXqK4gSYpSbs15wtDnYJ5lJCQ0cwdE4JFpx34q+m7yq0thai9U32myyAxBIS8az
gZL8tgaAOcjdcvY49afda+GNwhGRokq0En/V+FVWYAE5lWbH4Nnm9RQuqA/RzNM1HcxzUYT49tY+
1I228JBz++m8aQlB8k0IVurKYsZmmiFy2VK7K+tYZv2XXX7ZS74OgA90adzEOeFdWkPcAHnzTw6I
NhLvzule77vdxcS4Qqy5C2b5wDsPfCKDt8BDUV5FOFIIfZoE87pU9GAjIhR2qXOnft2UBMCjUPha
/235jaDfGQm0pLaIY8lbiaYBPwX0RXU+XozUnY2toCiVyJKom3hJasPuAHR9ThQxzK6XeYbG9OBl
s4U07Ru0DxufVyLxlab3Z/L7v0p5mFtcqxgpw/97/AkVq83I+Bx4sGPeDO2S8NAqaTZ81DVZNeQn
VhCcDHb8AE3fmqYoBbKxtLdwL7IEHYWz0rAogFAwLgRJ+Qyey41puJ6vb/plj+v8GZc5imu9OaZO
rw1Evdw8HxwIIdu2ODLD5ZdQdDUUnsnscizl/rtX2OtReQmXOuqQ7OfWVNCdTTJYlpRxrU6GRjcH
ltfegEcv7Y+69xEkdvzOQ1q1/aTX3i6WpXVs3crRsmNFrzgkIV6WTmMhtjx6mCVePl6UaKhLLdoe
sXHTo00hSCqUFhKrIjI0ZY5+BGtiEg57Ea9Lzyv7a7/oOyVpf4toJcV4FMrpiiI982LRJEZBVZCx
B875OFFJ649QHFwaskCR5XuzcbDxpfTKKodDaxZAcnNV6heud1lN5Qf3cR0uVvXLrScTCidNnTZF
r6tDsnuiOn5quaYpDtXN+Wr62aczyuioDg2OlKanW6WRSRVvZUnJVaIYiJw8UT5Q29dIiTccGyNJ
gbqQ/8kG1ZOauhjgnwBqXaiTfOBl/Teblto+t3maafCwGjp4R7Y26bFKn40CnDTL7FJPssOOiYjO
3REoHv6A3CuK+OO81aJVmDHsIn+A9R2nsfxoJFuQq4w5dD9Cs7qlULbGwKiIZuiVchpymLPk0Faa
DUrCBUvpUTPH3Lz5cZL9ITl+8ou348jwANxwvOOc1GNvd3F908a962/MykCrFfEckNInW2REXxW+
KeGNQzStyqtE3bjR1WYMwtc1urocXR0osBRpdPErUmigA5RbIkaOecsNiYFSYKawlIBc1LRPOWXN
7coXTTRdTxYPS/wbeWsZQ4t150GMNUhzsMvgZjzfbP0MGKAbj4pj9QWmWSidaJAqdJ/DecBpY+q5
3+gg4KAC7R+A8uCeAX9OXQF3RmIg2NQh+jnA4EBnBm8UkZZTv3kdB32ESvLALu/pBGw3vL/6W3f7
J36KvrQnOb5sA7qRQAYF3Xd/fXESCCtmT0CYxw5Grr7VZsT1++NmQ6rjnPULtXv4YhmbDv8XUS8d
Fn+db8eTtTE0/1rctxZ0FDAYObdwAo5ZWoctJpWF/AwRZzzE/NQd/X1JXiKvzPsRkY5WL8E6pmZB
mTj6kUz0nx6OZpwI9sRmv05r4Y2nIozs7P5fOEvWTYOMr9FWYZ+i9lRYfLHD8LPLjQAK9E3GuIUe
Rfiali65ZsFUfklXFMj6r93TGgzH74uazl+agDt+xN4x4YExKA2L4RdGYSZnBOymXn7lUWgadUhK
+GJPcZw2Ff6MgOZLTBjjUSdv0lWY7WDSFYqn8WQAwBI0q4CVXO1NhaDpVT5AqpM1LPofqjdQdpQu
wgWmiu8pu3BmtSMs9AdaBA1Z52JxR/YbpkS152DA40ZxvbsiZV3qCBCDQlvdbRjTRkG/0HDNa7DI
AX9c/76fxMRHO7HMFbYgWu/EhpSuI+v9IRdV7OUm9dvVgYCv98ODlxJQmDeXq/y0MY2ll+1n7FJs
rUh+SrVB6BevSeRmZdeLYVZ1xgSW5ys8c6hESi3tX5fKO9dzsEZYmfl+FZtruLsQ7Nl9godUFrf9
c44K8ZsRks2dQ3DKGwG8RdakUA1f2qZmk/JIsngz9ZW+GjCkfnKmeWcQDaC+K/jA1SRWyStykxp+
z9IOScnMRF+gj7ECMQVJMWYGuf8iWF771JHm88dfzpHhhMNFcA4TwfjdCNLyZaJeqIXM9bsP6ulO
XB/7cSaLOnSuzBYvBm1ZvbEL7LNFA+JBP4fgVVBN2FTUHXcN5ZtFNcr/YA6mvASnQIF8oau+z7cJ
Om8Ptfwk4XuBQVrnjsAUlRrYE2x7z2JpdWYtlu5hurcQPLeq/LKdqnE/YqIKc+OK0nhJh0/kTj00
R/v7dr5bBjy0m0sNM7qQdQSSEZC8Q1KrMEbOyp5Q7cyF9LhPVhbJQJ19zrQJm6u47taKhiAxPrIg
jinAwzqKyAyU7b4yWzfde4joL7FC7Xy/GOAvhIGh5wTH/uK3W6CLHHNSss8VCVv8J5gja2Erc5ri
N2Pgc/u4cYpMDm1FxCHQhuAUVi9Izc/MOd48Fcs+RqC5xMd2KKP2YKj37DrI519zY7kq5CBU2Vbd
wme1TjX2JSYwf9/Q8Evy4X8VNmfU1d4S2V4ZKf0GcBybLmKyNpsylRfFv1iTspJgtRJL3jlgoam7
0D3HCLLBe9rMU1jq82dm0psSYXBdJRad6oxkDWxlyWR9n34Z1REJL3JvOyq4Sp7S1Tg0GWbnFVmP
AdTtykYi7M1eJGTI66Y5gxtDMBHkbsS/y3ebblX5+SZkcqrTRHzITvdVWSpTAu2ZmHcCcwPZQ0vO
rF9UZWXN75h/FNrZwtmQprKcoEfOQ4mkEAGNwQ/QyMpLOoxVILNA9jk4EFuqVz6tcQM709+A5TJB
AYwZB6fkvgPRta+kaSbSXby38CWI9WGC+aWwqdqc2+jZPeec1aeSDv3fWfAmITDTG/CqizGuYgoG
9BKUfmGRa5jp3SX1Rhl9NAHTl9hhXF4iTA74u0jVj2hNC8cDDBxC2mOMgOwCyCezGqc71xuSdi+5
sYnojyNrkD0P64UQiRUELHtS88QQiFKHcLs7sFT5dclvTRjYf/Pn4p0Aq831ojmFJE02MsaL609M
nUh1oSeopGALMS1xOX0OdKgqj7qjMjf93lmZk80T0nomy1oPnMRhzS4Ly3wd/OeBm2HY2eEOztjX
z5L0y9NR0DZX5eIIIyzo/f4vDKhAZFkePcR2kpGPMG/e5TJOqepGPgWDyd8UG30opy5qoFM0v01g
klfiHl010k/2YL0uf6m4XFhYK7/tfXhO6otlvbO9nqPI2UHEFpNW4sTeUS1pdmucCvvwYW+9ldQX
5BdiBWn+x1lxAOUMgbs85fquHMUO0C2oYlwma+PALurQ759Xa6F7iC7ioxJIt2E6U8W7SE+qxTX8
8+0hT/4tP3XwGH3KV67xPyAvMm614/t29dflFsuQ+4FQkZpEZMwpoZXH2OiP91SnE3+W0AQx7Ahz
z0PetIcFU1UpL1zMfWNqbLnhEXKFVGgPxh91tsavPUYooJhx3z6kd6Kj0SU8HOtYhxqk8Pml9bff
7pLyhbVamJL7goVk/Y1YXmnqKbgTVF87jp+y7+TVcOZ/RiXJIPBEiA08mU3wzgjps85W10ST+UhL
ezTvTvH6HreTxr4m9a4yH1ZSFUt/conNCCTLryP7M+N7RIm04YTZTxxJImtvLu+UmCJRdsry/uPy
/KZ8LzyntOWxMRFO9JN3DOtljUOX9S0R3B5qEaTbT+tTpM+9AAg/+PKNQNh7ijgX2h/B2ZH3lUaE
IgJwPf6B9sXqCgCVn718KfzZfrNn6692J8BPuhEDIVD5y/iu7mzKbe98vEl5xOGtpdcXAYkiUpEX
Oia2HSzZrD0Nl6R4marukL93potj9G2fQRG7vX7RH/c4csE44ztOY+TOi2coTls8+56RKAZlla/s
kqqi1SPfmOrtjQ/CoyjPj10eDpj9bVmudr2qLY15KpJvs9EJj5YqV8vaIvxgG2IhKi6j99dgu0T6
YcEW62DpGw6BbEzIhSXWiPMT8ks4dVJaTCbMKmkAFBO5spLeaMmSrOQ9l6V7W+ie6vbwpByaJJ+G
NP/TNh2RtvpBWqVAuYhs/eoZxr/MzaMF0ed7EsYH+EN/witO+SWPjFRZsAJwLpJIYMrAbefwob2x
C4EsmFyaNAGjk4c2H49MOK9/UVyzR6Id/KI75ZdhTsgP0S/dYTU/5TcpWh0iVAAcOWsnm+Ick+1l
LSYp3SfeUnGkmO2e368AT9FtnBS0TdtGJS/vQNR26f+9F4JAXCSAnEYavStE28H2MCFO8MKwbuVx
ZX+PPsSgc83PxE8vJw/h2NufC382LDVM6Qfa7lSC6BENIWnEslPr2aEXj66iZfzS9Nd4T4+zMft5
eYApd7lajEXWKonaX+bnEiBNLrRmXPlL2gNpuX4qk6bO8x+Wgfs8VIWG7VBY6auAW6wyuDketyUI
ebgnSDv9qamBmyqsNP9g0YuLmu9QMXbJtt2NW83rliqbQmpgruSC9wxZqOzwO5DK8LxrET3K0143
u/AAeS7fQXVFb6ZVaDHBPA9NniipKEr30NgzQAylDt2/9Me8pIXXZ1briz6y3LfwX2iCUDoEXMV3
cMfSAcYgN4KQ1+OzEwRT2uGxVy+v3DJrMf6Ha9FnTp2AqrlGopx4Qm1dxxr9RNR56VnipZE+RdJ3
hXm8r2FYVW5s2nEr0nLumJh2JlfWBCYahgyYn+dOGnH8lnD69RrhJ5prunI5w/ZlkshuBQn1qNFc
6JAFv1HifJdSUEDImiM2CpXlmF1ojBYrJRvMhdcFH7DNJH1kFdUtwGWGLe7N/fwfejxKBOW7uxXL
w5PLntBqXGpkdSSNx+gQe7QMB2V3K12LiQUZqf5rU+9vrzfFNuF+N6CwyYuPrahvQP2QS0dBO2ze
f1hwgcXsk3HJ3jEisoKQtbTqaFu2IdeOvN0uIp1xuuVH5YVxowAIt3JySV1AxLDpgAy52JshGO9h
rpNDGNq0gl1lAn+hFYkLGbPhRbTQXrF8HiI4ufeFwMMshY3Twy1eFPH4DkCDoyLjLBIXYQl5jzTD
p7zaNRbIXfAhCx/QC2Wuu8NHVOo4MoFF+/E46OaWNMVhXnbH2nCQyUXsnnYc+3DLx1q4Axzjswpa
l/59i4SGTi+rvEc1KUvPwwFE/wK039vrVNu027SNZkixqmWsEvu/a/7LnquLkwaWZOpx+eVbCEhm
RxVQ5kUtXPQAgfU6IMbyqg+WjwahStc2BlrYbtMuWuImZtDteelTw+pO18WJfjLQe6QnDXdR5G+j
Uji40MUf6+mt/O69nTzapwWkixXLyQDR3gpBC8+o2OHAQ29piMmCGcgKlIt0ZJdVSE+3JDrBahWz
IlwY5fyY9/ibZltnhMNC+cqVe4VDBE/rNFuzXkOnk52Q57mw2a7wP03dgtqG9F4M3sFFnPmALHqt
Cu36ydpMNlaCnUmLJ6GjdaQ8gBrQHUgSHE22gmCmesihucBANgxHXY1JI7y5HY9HwKL41zXFqr2x
PpahgXqPNRXV1fqAojDw5sCRn8NXlVkE/IdTbA1W6iiZLh4gbPfIi8zcGlXgiQGxLUVsG+vVvh73
RD+s8io24IiU2UBTIz1EUvQJaC+KWONuPN5K4OVRGRVzQA2l6XDeyuto23z533iXhsQtUBwfEooC
tbOAhcSe9jR+1UsWmJ5ZPvXj/ijhALXF6iaem9wNB3A3zyyWXDdXQ4hHogmFwUNWWuGPoPBvncpl
mg/jzKM+4LEM4HXYH+BuUzrwfSMxpu5SPH6H0LrJfVlDikXyvD2uM38jN7rhRarkLAhfsF8Oqk7J
3LYz7UoWwUWwsJU2bE8+KKmAO8Rs/izMXn+0rsNCV1mCLBzR3++c7sz11zMytMfCD2ld1V8tGCFg
k+suEdm23oE/TTeKCXJ+VGHI4m6XfzlcrhzmDoy8e1Vb9Osh4unMtm2iFWbfW9cBE1pR58FgpE3q
o8XGp6h34ZtQ9zSSCwa2GBFl1K6xeKUIj9MFb5uWrZE40crN19cqAyiJ5BYYHpzuBkN57xW8RrtE
TKsI6W4MMOM684AIwJvy0Rhz0/5wlbW/wjYO7+aLC6f24arO74lh52mADGUcrikmNSnBgeN1Rtd7
HVFbanRWrV4A8kpSQsva/e6vrb6o4NJ2r2fbkzOprYhYf2aTLfZ7NIos0/fzlBPa6k+itCXBSfZg
vwP0R7ZpqqM/3JWUGFZUJh2X3mitUf9qDYd+W5DNWVmLSaINymxZ8WRSbssH1MnanXk0ypbvrByB
ryVcOYr1sk88pu1G3xCmdbxLrr1fNuLZoi9FhsTWrjgVloYFNwLWDuucEJ+KoLS1ozELuick+GAG
zjLOjkOjzEvD6a2jUunO032WSx1sMjksu9PSBIhB1uPMVZ+W0NHm4VU0M1EXHvM50oHONihr9E+X
s0DIPYbd2ZusSoxfxkuigvOD4hBO4FL9hB3Vg3Mh4xwkzTRCOGxlAFCos6nJKaAYsRdq43/RJ0aX
NRI4crxvfR9rg1LMG8GooLP6fcnomz1d9qMlonoV01ggiXu3bM59pExvpA712pImL3IEy5/A7M8R
lXm3ylc4Z44/If1+eqLCVDSs89lmgTmVedNRFahk77cheMxSv0UK/21o21RzlMT5VlqcvAOO1xq8
nnwoC1bzqmPNjTwgFt4ab5gAcK9PzFGcPZ0iBGMob3SdsYD0rgsuMLDQeTKdpPPSy45xFQTY2Dyy
4ZQzrTmZ5dcjul2tVtjPtPQLMoqKlpIWG8opTYDb2w/nWidlThvA4HY+oP7W4lyNEXQp2ga3za99
4oNYrLobA6avsRkUseNK4MxZYjmqfgxgUbwE1DvWLjWAmd2wCiL1W7MoCNo2vDfgqoYZey5iS2gi
coLj9qKRQWgTGbMeQws38jsbOBaqbMYabmqAVTRZsyyQ05A155IX0Pvsa3QvEb+JQp+f7n1+DNOm
TEZn2d97MOgEDuJd2Dx7/X/QevXbnIP2Rm9CM7u4KlLi4mDi3VMLeC1yn4EEKz9za75YV1IrgyU9
4HdMZxwIkLbD95vrD6pyaY/lUZIuzV/vGoDXJA9spFpAbhbWgPeCEpawtbN9eXokDFPrl8juZ7F6
hi2xfGZa1fYHIxrhXFzNhBwRWLxZbkMWjVIM7gfHRB9d//cVIwf4pZl8UNyXDSZRwD66/RjFEuw1
K1zfzhCcA7TVBVekkcJkjha2Rhu0SodGOn4dUbqR4fTGBq9/KiYYSelT8E4JO5bbKJoWKv17BSHF
c7DQqSyLxyqqLaCin9SnxOOZAOsx4/H42aGpUNSNBfxka5Eh5tKM+cuaoCyCtC38O5JJuzFzEVGa
5O3HL4uQJ+74sRC+5ELIuoSH08drbXQt1CJuiZVkQWtojQp3XoZdURRR/CvyA5ZSeMlS74Z2S+dh
4r8n+peUUrN2xCRapKON6DpWPmVrH8bsemz/PVwUGisKtMGNh0RcRl52D+v4KsGCgr294zrE7H+5
0aTgciohNjWjMEi2RAu48ZrWQKIDbnx1YPGvEPp1hs3Ap6bHO6BIhxUmtEKAVrlS7N6xXfUPtwgI
3xuS2m2eh/GpZXTAjUPtoJeF4Ewbkcv7KLZqyqsuL6A270RoNwwCK8VL95mGtUDhbCYsAFdblWiQ
R1UjyjFZSDMWILQS8ipezgOYG53SUbVEu1bB+RTfH2GLGzG3X+afdBdxQgXrP49Po9qWzLGRYV9G
M8E9If+CDRZzYNCUNmAfl8yoxfqbRXKVetqJZE65iJHdyOivFboBJhT6R48nsoTJL3envlbAYecW
m+2l8V6qhjHp+jhZHou8Cidh5tG/frXaA5yAiLyNiPZAhhPnohFeFcCGUG0zbUNuXp0BCopnTtuH
lYB7eXXXwvc/T8Zbt4Fo/yBxoufoI1BJBHdHmQxgNeKPD38/eE7kl6phSvBdAdN29qhFQsHLY2/L
R5kpM0qC9oMdCNK4wAHUxA+zAhvS1KrTpdKUAy2Ho4zP5aBcPjSfyYgoXd52Vgjb6KgFMidYBoAS
FtOI96Aj/57VsndU6E9d78lgnlOkUOeU+WdhYoMako7ISiUUEGGXD4fX28nNJoXbk0EShibHoNFv
EdAQnT2bFKn8m9ycMRVzFSYnKaGjBSFFbm+uPVjrCCbwU/H/GnGOXDH2NSDqg7GkJ3NboKs335gU
ZiMTZ+u0MFBQ5XBDv/t+VYIITYgCxXMJilncgp1BOFi1ToecZ/2awapDGYBze7JWxObgq3iTQlHD
KWw2izgZePp0BskBCuoRPL3EpP9Bymmm1b6cjma1ZXMGoEEdFle6mn5jTbV2cQdm1/f59FyZAf/8
JkuxoO3SEIYR5bGguP8OOONW54LnrsepFaYytIEgjRSn6Bvsk51sbXWoIxflZvsuaSUcY9qw3ciU
pkgm1pAdW7O/LXy4GBkl3q7aEnlC02QTkWhLyXr5ahgXoZrPdf3pZP7+dk2b8igL5LT35FFvL5Rx
bnuJZRs3E1JNvEz2d4j4XwLgkwtrVjMfUKACRBVqNWkPT8fQezOIW+jak3wMhiQy0LG42lAUmvCT
1JKJC0azXUjpDM7rlwZjVG9snlpc80q+X1lNBxT7CmSEmAtkFjuY3cGsMqCcsEuAxlAPtWE8DCnT
Q2btrhDaC9CvkdbtmNimWGAIK0cJcfqKZ8r+sPQ/fMaFhsMwaYWxcDRfdx2fun4J22FO5DtNH9sK
leDoj4J9GOy/LXPeVD29PUhxkernQ8Qo85EzdljglBXGoId7TLzlbmhyHeLCvWpcKpxQt9d5LRum
HkcQMEbY5vifwcuv35f/3yE++Aqd46u06+T7X63mFRJuRlC6vhaCyUNkQNqZPu9dB2wDyv7vUlYk
VBS8H8xh73gOupmUmn+p8urf6k8VhmxPvE8VzmRXt5P80eF9JzfPHC1aQ8BHwn/2rzDVAHrBKz7J
v0qAdFHvEKP9YSkBdmdt9YjqwYY1VTf+vTV8GT1f5RzG4wxtta1/b7z1A4TbQtrG1vdzrcsCY8Li
84fdSinZZBK0FFEMWZ2eCCjdgKkWXLqJMlarIGlFUPqdKmQzdNu87mJ3hdQxgTFW+loIVViDHhix
JzhC3mSMVO4k+G0xZsdEyZJx55svJX+7D0MvcksEivYk9Wih3gS4aS5NP3SjgxdW6tK0wW/Zh5rE
85LL7e97c+j46MXseu3VaMveL4iHY3EEZCTRDtcyP7+qGFkEVz/7sB+0m2kDwh2CgCxophmw3r+a
WKVCfDW+8zSbpzksZCTtvtwYOsOawv2n+nw0jvEe5OZISdT5TgMqTWDbGG4snW34CGwZgqJ0WDPj
va5mGcUCkjuvOXJaNbkhqKnS5rEuak6xQkgBHol54PBEt8oFsv2cipL9NwN5SFb0NXv1O5F1XND/
6V0U/KFMBavJtIyr5c3gOHnqh1jUCjzFEW49dt4bPGadqkOJXA6n3c0WecllKo3ZCPv52bu6Dpwb
0anyhCGzbVsNWupskkRlWD2eLUmvXpETQLOmsrGB/Ljy5uia7yw+UD2ZNaYCgr5GHXUmUDs7Mcbj
rW+AvzwxupdaXwC2sEK1hEQM2YEBk4V1aGhGWYIOq76d16Ao6tKJpBhPe6p5NW3hnaqWO2t5bpCk
wLn9oLo0uhw3SHDpNNJyappX27q9xJsbBy3EwOEDZC0V6z0JYBKesXJ2aBNPNr/ugBnu50xj8qTZ
dK5AzhxLzWNsaa+auV8vKuNQuR407KKwwtJxNgCvL/TPyAe2Kr5LbYO72g7PaxMrNiAFwhBd/yjH
IXn/+6LS0lLNiyKf3qa1QtgNQi+0LDrwXo0Ut1VLfXQpkz2UTsaPOzWj3XECLn53uQ0D9e/KAH/H
kDHScigI9H48J0i0W3l5g81ExbfV4sipYEtB72s0Cl2HI/qZWYxD56dqL6VcC8isbWZiq04HIWhW
2re4zrvEoB8NtJmRzWRBSm3HGfocA6XSKCWruvUuDoSFsqn22v/WxbZdkUFPQ0riDkpXn/0Bfy4y
AQ4//aiLfjrssKR3o8+nhQci8KD4XClOT373raHwTlNtKW+GiGiw88wYWoMhddHS3V9E/NuOmXTD
IJmoqFkz5kIsgt6qWVp51FyVm9tIWRW+RC/3qqdiC24JhvEH89JhfpJbk56ng1vSY0DfzcG4/AHy
/7K4RVNjpbMlTLEF0L76yMYtBCIF1p6WdvhwYrln6c79+HIzIfNzcqW8Tm65LAVgX8OFKjtnJGFS
KrDRXVj9IorZfe7rDvynD9zQ4s4chibw9IZsdNV0VHFohDrx7d60AzcLWYW64kIhzDsiF9Wv4gI/
DoUbYFG4MXCS0WCPfWzjrWSuJr5U0iydy6Hv2EY+MfD+j6bAotZ1h6JCMXdFwUIxVXiBC+d3g6v3
4umY5n9RbctBIY+Vxg8vlgpTZ6JLmdMucRM9WQYfhJLElWod8EeKgizvMY9YzRV47H+wMhmywjqJ
8iObTDiq9sPDoI2AWuj+i0+EtRy5tXb7YgIEIGZzJhBySwSiS57WJUXiA1nrf/JPc6kJVCilgaas
i4zKtqyQs2JN68dsNi+6gDe3WN+tBwuLVTW7feWi4YrQql0JvfcndxJSlD424nqfyGdEO4PqBdmV
WtRYDXTl5UozGMZTswnsF4J1gCAOp0vy6X42tKWFRG6kSPJo6oVTzEQi9aLBf2CszF7lU0pW5oyN
vOitWaQEUcsNIEh7p7ctfyKp/yT4vnAvehnQUdc+BXb0gh/QdAwgWRq4+GmW+B8RtvHFvJ4FK4fx
2dXgGDBDUWJ4Tr+pSKxffWik+G3Lj37mwdrjkALHdgsYTkeofnrdwoJeabQfb2iPPvMoCojU5bpJ
wZtzoj9yavj99LDp2HYbf/iogkgWN0EEgz5aEWTXBWpA4TDVPOCdZ6hG8zdY9cAmtAIk/7ceLa+r
FL93NRwrJCSVVOxBaOMGwZhjG9EHMeM8iJZMwTpDHb8+iPeRGI1/wJ4mMtJKkdz/vZ/ZlS+xwzsn
V+1fgxgHRBSOle5mpt6FURAnTZ6M6gLkAHfjLPDbAxXCDGBoDYtg95UpJkiimn2ejCqrLV7X/wEQ
SV8PoGyzm/Hbx/v2jx52Jq+AW9PTtom51Mbfgytz6zO4vQLjVhuww1zF7l15ZzKPVN6KpI56tl9R
WwnxUv6IFi+baMgOJot2eOZLLPOmfIq1GaW5fg4NfW3oc9pJb193YvcwCyp9WYZfPgVZjxoR6RfV
NUgCr0SqjoG3yXWulR1PAPfcA839o/CclUweZrn+b2IycnxNzri4NyVFseOOzl11gdtlE1SJofXR
lGNiGnrzDBp+xhpTPaidoPyKXsYuGPFp0/T6iWnyPAmRame/Iw5nt6A8n0BsqMGjKBOP72uzsecX
jo0ewSzP9z+4JQ9eMhU97wt43NMdEAhurc0wcmCLj1mtM/JQfeJhDXy4U2A8ki66E6+o/lx9zSaP
l1Ou6dp2n6dynkM2Atx44pwUuwsbs9SabHqAaHb2MdyePFvHOgnBDcUtlcF9tOGx5aCsHjy/9fIZ
BHDJEtz/4dFAVo2Y+T65Uu5y31+LeMU0H2Lrgg0sfVG3DbN/sqAWUQ6wwyD7KCl3oZeqnnUQFGAn
oUHiIBvubfeL9ubwSFDb5VJSZxUgX3MDLTcJFQwpddy+DrES3hbhELZv8iPAk5oK2uMgIIfQHVrt
kL0x2VU+SI15oJovCk4pEtOcNAdIfmYUIXOirc+JeS1OBVo2m5NuMw3uhiQl6/FGPUIAFcWPeYdl
44DrbSYQYmzPh0k/NP8ftlr5iok5FK7EyThpu+PklADM4vbYGVjqxPq1b58gaWYnBPBe61vOhehC
pBNBP70m7AB2ExEFzzbyx7hVfa2l0d3cTENA4Luj9oySu6+OVnCGmptkcn8J8T+qFMoHccmPIyE8
eZZ/blg2yIBWSgTIVYxZQjoZz9xQHGvJAhBr2Gv0Hgs2bk3FQmweFmzLbjrN/9tD2kxtOKXDW0tE
kGvPxTUIGGWiXXWeMEpRA/vIuvHfOUiD52nkkH7H/7UUM5oR2lGFdW6iTjTsW+02WN9y+iY57Xju
pSfCe8dUngfwepoIOWB5Wy+OHQ+D+uaOsCzMEmJUt/1ThYFsdZq2nzNBrLY2o6usJ2yNCEW8hr8T
n2McOG58Sha2fLXXpYtdRrTu4NS3Eqj8tJQ6IprslhD1V1rnKiNVi26Ep8Zl1hRZ5HouzRVwBg1X
ngZuoGBXGsZ7stk0ncSbtQqbq2kdz5MdQmh4QsgHN8kblFR+WqxJTqp0aMvBQn3PYjVWhgCm7cFz
Kolz+XEdWg94TGAKWEQfS3EFB333zfDCB3aBaw2Ez3tCSFNq4nLEGG6p14JB7OytlUdUHPYUjBAB
eGGRjmjAVMTJDEWQ1/w51QHQKqPb7ZibSn194IMXC7E1g+hsBAtEXzNwKKcMjh5uInmxC9D2GhOg
LQNG0HJvCwYSeVRKewR2pG8os2flLh2Up7ZjE2DC/q51r3UV6rjxd/f3UGfp+yUnwYd1KWQbfxCo
oLx5EdaghWhR0Wd58D/+VEIw+hQz2WmRH+d6iWEGDqYstCtdW1o76YHea4XEbaaa+gDJHKmu0tc/
4YOUbelnObIyblcfBkMDXDPi0kPFbckRIoV0FS3cJ+Ih4AdDwM4vXCKQXzDe+Fxv1UnpciLox0S2
Vxnj4wLE+fqVOlbQNtxUb0sTZpma2SA8mp9mfVOcX0+A0oMMyPC/DBmGc5GkYn47mkm79k+g4Ahl
5ChqLpiPmIwN0CgD9QgSj+/NfmVfGFNBVrhpX74Z+KttAkgMm7/8YuP3OzHAwT5Fi5Zmkmb6fkry
wrybRChMWMWQFVl/OSgBAma14OkuZKfGVrYNyaJj+7neZ2GzyTR1wGaCJC/tBfG0YxWuzh2M7V3x
uLKrNld3381fr9mRcFRoQTOB+1tStRXSQs0158afT6hKfWFe9+dXL3lNZYwdSPJaU7nM6+LS9Ipk
9WN1W+phNK+vkIyn/dr15ooA3nMdPzIOSB07iK5usKTvRDhnvDs+/QrxpP61qwe9xOlzjriHdePM
7tPwxv1bVOFgFf8xookkOSIjZIgPfZ0jUek93BXmfK8T4itQAq7ONLdjEjQUdqsjgwdKpOJZA4S6
5xz+vFP183HbOJUDHdmRlm5dkd9Fb4zNtpO9MNcV9a4//ku6n7Q0BsLLBs5lg1+cmbFdFihSDY6p
NmDpmKpK5YNml75gKKLMt1z06p+fIyjHofqbHSeQR42WwAi70dE2kjLbTbqMdTPNggRuZG2T0eEz
An3s9S4GhZ6IrV22WchoE3Zkb+M4Zof7p0K+1DnWDyZ2JqdGl0WhUxHE6h4WIEnGPhc0KhoX4SyY
d4t5ZMl1cgkZuhC+18Y/FoNwn5NvamK2cuB4PsjgOyrkhHKH65YQkTm/eUcYSDNLUPsEU4ACyrzH
hDE/oZaiGTpw9/50G37qR630uvBOtsSoL2twrbV76kQ34XMfaCYkJK2N6HfCxt1lS0BCpdQw0uNM
Af47y2HhluPNPdxvvbKTkjxuibcD1AccCxX6oyy7PqZEGOItp0ePbfFDnmvAsU1HSrErikhykaFQ
GO8qxoDR/hncckRRR07QJQu7P09+ENsOKCi8Nf3nYma3s77BWGkYl5mTglI5JxuxpJbspU+Kjv0B
7Q8QZ7DOSjmYAfT6Ckkn6QoSL4fY7hSy375EsXpuyzeht6uDTf9cIYSI362b98e/CTyx+mRf0NQ6
VP6WgfbP2cAxqNT7RuGQCIl19XM37tkcB2u5lLKaJGRUEOhfSvDieREsX+y06pBNBPkbd4qcQbz9
bMjJd8NU7hS5j56+zQUutE4r0jnozM1CZIiIwxDLBxw32LlncBN9JHRzDxRzFg6TzRxxskqNH5Ha
X0QK61sy2Fux51amIkexK3qsYldiFJKEW5NlsNnUxcyI+x+pdyk3sbQEKDDZtY5JWKcfJDbKWs6t
saf0/ONnFgV1Hb64SaTmJPrrKAXTJkkNEZ0sjGAArOuf5pqoek6uV/Yr91MGXnu+wvPsiKxjwH6Z
syHmBeIPDU8eAD7PiqhFT1rOb0Hj/UvvHAslXKfbRF1OTFR0AjgBiTdQ7BhvfD2Mofefgjr2k7aY
N/s3SDYYeYbw0slldSBBmEqtW4mdakxoGHNRETKaBQvMX+3EaRjOqlBOrKOMwqbGxFVrz/IPCbLh
L7abu+bUIwlpRqtpNcchWUaRZ9RaebLQ3CP+ug3n2c1uJhGziXowRyBzo8SXWnD93BbCxI82nzRf
cGN+8MptqPR8wSZK1hygs1UcgqDZAbNrpYhxhvFqd7fN7FooXTHDPGF+uHtDFQOHGdmCuCPJ1nPJ
ouD6j72TOFs/4Ru8uvTyTj5+YzIgJzhkruG1CvFENqY6ku+vu8TZi87NNDVZRtB3u6eJwEBZAcgE
ocn3tWLqyqFacmnDR3uNAMY3oUFgH1e1ZNx/R6NiqGCm+kzwWJGLHLipv/zNlFMFQOJFVrRXXodQ
fkZ3wWyf7XHTme/7Zhbv3st7WtE73uPkevfwFvXM9rExg0R53HUVXIN63XSV1JEt/Np/s1J6TqkR
NAjwCMGXxT7BzbXbGjXWpBvVnCiP3lEhBBtRfYQgGggNsmEXVYTUUQxQBTnNBV/6NUMLdHP8WEzW
vNRubBb7duOWroktIN2MvK1Xpfbk0aFHe6Iatc7cBr67TnqsH38+8OvRrB6bbTcwFE/x9qx0nbcj
EavPvLhmrEFNOAZ1R/VSXN6jtAKyEfYs0ZSY+6x3NFZelNGU9e5/v5BAJEhP5w4Um4T4Nf6SGQDo
U//O5u4nw56Q65hyA5Hhcnhn3GjWYan2bSHvDhP3T4RsUU7EEtKERh6kWdZh70Wwl9GtK0mKVlLN
TfjII1h69Jk3gnkrpc/2fP7TAyCh0wcSZSscID6vwX3WN5n/cG0xa3UVYEhwJq36VosZ5oA6H7Ku
KYqs/2bXNbpGt7N7/nYp2deKRbKfk5wdQa5qBnHciQrqnsBp1S6XurZ3Mlt7d5hsx/MH/t/Fevtp
AAJ79NpLgis6kOgaAK+27Ksv7ugoqa548A31Db25GpZquToHNt+5i5YbSiMYlpqzEJyDod5Nq5tG
RGz1gYn6VPdFY8bQMdA/USYZLrBUr2H8xZUBmkpMsldkzhZFqFfVhJW3CUtL/hueDVrHg6pI31vi
5yvWc8U85zRpA01TVly0fjsmMrReR8+LKOgq1QGgkYdOAMqjFLyOvHRkThEWVbj4MfD8AXWtJwpN
78FaLxbLb1KKpNv+fjQLgOlr7gx6Kzk9WgresQSOHHTEkHWU534YTTyOlnP9ogkOxkEiRQQZt1m7
mMBI84uNTOvUWGIVbi9lqqyYDfuqw8okh4O17fz6904Bpubjz8tZlT7xIVpSQ6SkQIoA8kqqlGy5
X0hLXTIGQsV7aajh66KfLkB2Q0VpNZ5jPQAQy5F3zHh6uJS8XWUfGBNxpDvLiHFT+ru31oQtsqXO
ZLbQM4b9xmF21n5OEenrVhG6YiQOX2OSItXSW7zddaADZ2MxcYujDTaWv2GCMYP/HC0/fL0d/ff1
5PUDK3jUY4x+mVJqOI8qsOwp1K9H8cxl4vOtdg7QZ3/7y8o30XLHcIay+iREDBtPvMy1lORD968K
QuxataN9uRHkKaj77Pv7m+7MWF9nnBMF9qt0Nok6d1qdhGlkPnWgcVxA8cWruWLqGuEZg5KhZH0/
TYv7hLCtiR+YwZ4r3zZyJLSP2yMIa8TVg7YW/kcUC4dUbFN+vb09GdCOysHfPw+Ay25rwdqDGZjq
oDBZd0+A3t5iNKA3XQQ6rgiz3SCuULjZUKgwA7WZx5jug1GEDhUvgg8jpaoSOnWpJkKsDO3/7uqN
7coCEmKwxBq92w2z2jnVMNiu4I0E1aJQZS0f8MS/ogTRvu/G2N3k6Yku5A2FH7OkCcvgBlruYXpS
nRuqWL7GSgH07UPjAmVUGLD5uEe8kYroNcucUSNMMaXyypgyMzHpVt3Qqseg0+u67lMsw6sra+wx
V5GUx7OfRSLanWe1lPieqEUixcY7yGSkl7A6af2rDhgCawrGRzxkKOIOzNXoSIKCjX7tVm3X8j10
mk44Wab16tFqKlsgyksKVCtTEqeAzwfcay2tg/i6kL2ZxkaY9wmpEPahcBtclvSiYjGba5PPGNhA
5cAzQ+nlZktrE3yqy2uJofb3ClGB02j7pivETyvJb7ZnbR6EO1bqEDYjB2a1Gp9P+VcVOt9IdsbO
1OQPKUF3kbcr7oLPWo3I9FqKwfpqktUoxClYxPH47XphGL8rH4hUwg9A0urvL61191vCB+DY7R5K
uAM7bes4/wAmBs7eGPgDDOVLidKv3StyqOZrJdh26Sn/qBe6Y7MMR/XprPbzs0fV0CZif+Mb9T2C
aWzbT5tmIkuEB/3m1sIjAMto35HoVAIAwOMJDyx291FoywiN0BVDOmzLTItIT5JQpRSdwwh0iFrw
pH0+KObttjtABFMzTHb7H1W34cJ6gHPRS+SPaVtpPEL9LcN14xzS0MMkDqBWv1l8TBuyuo63z6K3
nLseDQHOSYaFPmjKBESTJfwug+PgatL4qVx3nMXQmthLDtxZe9BNcll2AOkKA+6jRaP0SkhvEt0B
jLuc+yNoIQ0eWdpGDtLfB64eSTh6uPheWaI2IXF3HUEAV2Zg7KjflX9KXCBqcTb9gFe4Seh/FXYj
HG1L8c26LIvgNr3a78dvO57UByaomJoMGz/C7EOCfD208di/5Dg20fCdR6nv4sxvDc4Bygzej8Gx
a3Zc0sj10eYm6Y4BaYbRRO3i90Kit7TxMJK+zdeXGV8AqzN9xiB2qwShYpi1y45rj9n/ZhEtJ+z6
zfZRVp4dCQhp0MtbouZI60WsXxSvfahIMD2i+12aUW5TgXr6tHguY6YKRXorXyaPB1s40OKqOwJN
KKEnu/DKEi64tKa/J3I3dIfmpCizU2vf79I52faCVGfKl4iHztD13PvxnnRo3dLA2VjCpm3KhMYl
/hOTHMr5NQgcWJstbynyP9v6fxGV9VNlUHX9+Oa/KGF1GkCdIwuN+fw891IZeHG0bY7EOAnXj9Be
k1WvM7wnABATkeB6MxHm7AxaYAgXSSj86QGIo6oHS49AxBCUeAmrsKB6kPqupotFKJjbs1u4/0OW
+WcHkbwKIe4gCJ7B8HmQ1Nkg7J2vZ76OREbnnCLXjF3BuU8uwQ8t7zrFrP6TnSE9vEVjl+Q2BiS3
TYDUHwtAC7rffu6llfTTW7lcKgBYPISrQGSH7424M/AOBtCi9KVkRnEJ+RBufiOuXWMbXzpNSK7x
fryRqBObVxxJdSu2x3ynSICiIQ4O0vudkAa49hyIxVm/KnRyIR9OIYQ9+krTP/98nik0zIzknKAs
mDu63nK1yKMqR0nB14pWCgbbyu/Libw3GcEW/EabHmRH3fC50fQHEBfUUZYxoB0Z5OTz7ycZkqEx
jy5GgO80M7BcUzFayLl10Pn+dL2MxwWyPPMrEzuZaTVxCXGZgOfwhGpORj81Ga8AiQBxwLJI62sJ
4AHZQTn9eFO/3F12g4g0owchHUmLmDXVAYXz8MoHBvfkjWj4DIP+xGp75xQ/2UwcVjvL0sBkjozo
TIc9P3RoTdUDMdProPLjCy5IiqJfrumh4RV/2fWt/rIGTeHwVLlMqcV/MJjsBXrCXP5qSiJibhk3
cgJZz6nmhDBKUjL0/DuzgFJyK2kQtjAfO8iy78io7bL+lVfImBEWWknaoeBr/IaBhGwasEYFipbq
EZMTDTTHqB9suTXJGguItFO0uASpBy9bS5naZ+oJtQktmFcXiWtGILZxRNh1alAoQghbIUlMEZ2+
0qAdX6PFdNwDzmd83u+R18RnjNF4wafu9e6SeypN3VMs/JRAI0cLGrctYhbvX2k1FQ+XIxKbDVZP
zS1E7HMEw3byH7L4mm97EUKDBhHMchIdCL28dUAVpAr/keZLpeS48XrY3S9HOkpOaQ+7Qd6WxaTE
y2KtylSpeVkoDk0B0wkINYnoTPHDw5mCa4iNdHNUNnuMTCNYHHr0geMd8fY+7c2dV9z482nydLGu
iRTjnKCISpT1g4F6eELbu4PPZvV+G5coVG/3X1HEy18fpisIHh6mIjZlZaQNyW0XbsRMnlEZTfKk
yYGtigMJHP8oM4u4DSICTtbZhwCmFFm9tMe0Mn+Rt83zovmwyBZ2of+CX9igI+sIqE5UKRF4Apwm
9pxiNUk01dW7Eaj/frkbMIVWMx+eBEzplvZ9cwpVbSlQh3WjJRUED1tovwOKN23Dui3op9Yl1zIJ
zH+rUmIeJJ2bPu4XJcOQLcMeMpwzU8moO2kQVFshgqWYWxa87RtqR9owp3Ii1YRt33Cv11POdBAV
AI+derEtNUUmvKuXRUcSIjPpdk+4v9TY5gyhXdS9sIJp27PiZme2HbjQWtlUBzjL/FDIT8+VRYbb
dJF892rI2R+T01M/fZKyiG1Cd3zgcW58M0rAEL63LQilHapED86lW1ie9SalJ+u265CYYNtllysG
5wA3bzWJbIzCG4eF4I4gnOg0pVfxmdk8HJ5yWzvHMjlyoWpU+UAc+Rs2T5iniq3hnonjC6x8NGDW
UPG2muerYbU+yU4AubHJRzy5SPGZzscVXzFnNzghBiUn75e8jZdqNsxkrgIPGjG0svBV17KT+BpU
QPkKV+PsfNb5chdlbufCdpGVjV4AictIU1m8u8D4kizpRicgoqJLLCwvj98iQWWFSZw/1TQVNd+R
nNiPZgEl4wqsXAxYa4GFt+pygVK/3cV8/pROZWxeiWcbe/WVL4cMEUBFtHv5Mqrm9avTiYDxZs3c
9y8STqUA7ew6w/GqQNIFC/7PDpY7ORkp/jwloXwW3X4duTLAG3bSsAa0bMQ4h1/dciaYgrwLeTTi
QkK03Ju07oLlQu7cd1+9kNzPTA4yvw6/+UIrr8dtlWsuIvmY23KKGfozg5MPvcRtVXMExshs+754
myvPu7/DGSmCHw2RGlPP1Otwx1VXKPQdhC+am9cHGRgDWuerGhRVg7FV8oY9BJ581a3L0fnb+Q5O
267ZaI971lWyiFDMIhACOM7LdhkSuoMQM1G+ejo6nbu61vjuIouDASSrCR6vxePlgrPkPDoMHGj3
EwexxqmN/2rP2ARQ2+cyGIT4i3mk5qf9oZtPb36y++SbTbio3Lz3Mf5jOhRwXSfhsy8jmf/vv3M9
MPsGjV9YH9erxGr/0sJlWFcyomhMTNf6T/YaWDzGeZejIc72p+lzo2XWs9AsyJvO530QY7DZojWi
XMW0NhEBya9TundqGRKgvcjj7N+a37i8SdFK5B+q4Avc02WO9GfJEJsZ+HPSroavomsX8lN+MtTb
4YMbozqTtrUzEDpH41VtDfWyKuTZTk2KTVNL6uUK9+GLfcK01ijJI1W8Fg/L36hjcq7gO5qqDwES
dmb2TwoJon/FkPZn/N33uDeJbloDhqau0PnYdYxrAA89sZzXsYfv1pF7meyg9T/yUmFou1ZW5r6/
WSwz1VZ6oi2/H4MvTGOH0744j/PMutHpHlmhN9bsvK1MfA8/6XZC16UgfusNO3hi+qrOCc5lGlbW
eqeviC4PLkeQpyx70F/aAenyHdIxZH1njM7K026DTi732hURqvrZs4UY4dFgDGLEry1n4G0iZQXt
s4UzCkL+oqDnMSqc9khri0jRPF8WuatTLano0JT3lcsi+i6Ck7uMicwckd48IKVASvw3avOxNm0T
QQIZE861Hb5WtFjIt3qn0E/9yzqo9xMZMmlD7XgEGOVdTH3ip1etPThY1KjwnLxO6zAUnjnivuas
ZqZSmHUNjSaQyaS0Z0yEHvQw3fYUVqPHwjt31Ayp2AaZF19D4xL380bC/iDUOhw9oQ9jORx61Tgx
T6Bv2L/OeB3oto/y4iev4K5I0cgPMJVabGM/mbIR9EHc6LGRlC8WP5B4XEFR5qUujwkVTlYgnTDV
uQ03z693SRTKAO3970CYoLQgXiItfwIqlpH+l3vQ4qQJwrPwz9vTw7dpffMadSIJ5zwGGybNYg47
VmZGtMEANpNELefonNcL967E/ORk3SujJSEg5Q1hlVGK1g2XXebNlQTA9lzWqBRLgGebv0EbtFRQ
EmMMJLiGUDJmpwZEVwZzS+LQOYHsAhEI+c82vSByYYTDjaNx7p+n7k2SbHhnfcbc825ajAEuLopJ
yFpsfw+AHTA/p16FZpGbQ7qjrJPt5Rdsaww1F4TBuceRIWT0nmv9/aEU1hmPhvsboHbjAB7Yy/T2
LBnVB7WE1EJzSWHRdXVhLIykbpXQnIlYOQIOBvBUA3/W4Wk+EDVK6HqcojvXJq5JZEh6XQdKIdLR
/PY++njnDBqPPdM+mtjxQnLzHGp4M+xQwHz8VpRlErNlOvRSUwNE8e3PjYfTE/ohOfo3ULhIIhvM
2bEkHcuQW91zMnaTbeZojKFb2HmgUzQ1UiNqZPD9rb1R3pOEzhoIvFgMm5ccvhrGFhkiWf91+8MC
zIZVPHTD8FX86ZSIWE8ghb0BSoOuTnOT0SlwbU6Y3a1CoEKQB3n97akN+XIPciPpt876kXXjQE9V
AEKicxmy2/z498WMgnV4WQx/gEVoujUP0NfxQAucZsb1diYM0A2cDJVe0LnDgNGy8j9zlfTbkxSP
hjhbaXqWMwsjhKOYXv1TsbeUMEn+FenSEWMqT+AIl/jOtn0iPiUy+sRaTfkh0gcLDnsLmejQ5LOe
aU3lnQK0FQIFvlS05wcV3FfthBPQXfarEleLFJ86rKN4ocoAcbiY8HSGKd2EX4EVLCd8Me1ZEPdv
w5U4OD0UfjJueKMx+P7aX56l4XFBZ+m4vNCffOVddvtJyeZxMbtyJH8MWtPT5CPK2kxDV0hehwPd
Gm9PaUtF8ftvQGMu2BKfHrJlTkyhN8WvpFTdDA8wIjxnzRZYdW1/WpBaDhGlh239c+KfGSPQUaH1
XpBKyYBm0L20SCBxVQIpugvZZz4H3+v95oNyd0ks4K1GnKi/XHFWZqv5H5CZhZUXwWlShgiKaEbY
GoynVPCuQnINhyK9z+Wa9b0as6b3zOChPg2sO8HBTgcBUR6M61UrCbQRWzNybym+0X3ptI1C3h9k
q7iHS9M/0Se61q8YgzsuXfaldO58Mb+fS8YufnSNeg0q5yJ4fcFbuU+3nRpyknXRzM/rRWtj3G21
GV7B6POCBB4iMCdyOAdEZWTHrbk6cmGKvnsMmYTAEB5hnp/Y/RZtpOIsmZQpVST8eBUdM0phnLqL
RNOCJVNWXsLT9OnwNIFjpujSAlCC9wniI2uF7DX7/EKWudSioSulEZfFMaV0G20AWBuGj7jlvfmP
o+ohCVKNaC+drXrogjtym7dHvReyofDQsxqnjBpMwhFyw166HleB0PypZu9rlIuH5nXwieHdT7tx
h1GDyqoBnEtCPqpfdKm+3GODoW3X+8QW8YMLZewyXCBwooL64mptuScrV/WmPkNtCJ6JkLDpdCXQ
rzfGwQ+Dtu2P1jqz1ifbT8wA06spZeXt78/JYm2OpOB5GeKla/k25N1xppwvAFrr5j7cG1BRmWVM
O503inGaEeU+cDp47N6Zj0owq6ptdHR9FXATaj8214hYEZbpuq6x+xqO7z0kaCddOWkPufFAsOIz
vf48LHJCNdlGoOK24Ze6Sfl6qRdIhdKPxPTrBrQh1xGHTXM046zmKJm0XdRZmS5bALQekmmk8wHc
5gpYjLJEjuB0SZgDw7gjqYFqlbHSaUpxOkBpkaMYLJiqnq9FZinZjUCSGe1xMVGP2CZsKwvRKoaa
TixRJMK7nfEfGOI5XJeIscHkJNPZhRqio/6WOizz16tU0fGvrH0SCrWhNU/TUUe58K0ZGwbb5hMI
ftl3vvVIVS46ezf43NKEOJNHRTeX36NZQxG7mrzz68tqr0czq0rmaYZTydziZvIyug6oXuAKRMD/
gm4AXeedh9Yk3uH1ljafzIEEdAvwpGuFY/soAR0/J784Ve7xSb9hDffLBpijJx3KHMinRxEJ/7+r
5DoWSSrLqNOCSA83GIMaF3fKXm3lPRY01CwBqYJxrq5wO3a2xM7L5GpHD9/fn5c7tsfuGCApshg5
q8cJ4T8mJ8xXhwhbNiY+E9Z8Z47ocZmYJHB9OTnAYSx00t5n4kILbUigqUIRUo+guDr4nnfHRMEj
gtfSE4DBfam0Xr9rxAQJeY4njJZalDWiRPIoYVyX7oMclbbU+oJYY3YroXsSil/tUHwEtKC+2oDC
458ha6QckqEFGVqmh/kkh5hnRlbPMMoNmsk7pnFjkADuXwNus6hsEP9o40tYR+DY4gODjq7Cvhnu
FFEAu9cFwBzQ2LtS0x+6YLPovd8SWwnTKM+LBFE3dJMmfzofr/jBDZe0QIp1wXNfG2Y7Vyz9x3O+
VrcaFtFgjoeEkCyHtcwM5q3lZVAbs/4dA8JL72iHoLCsSA7iPJLor2Red+oAiwsgEvQ+bj5JETPO
w5kixFacXkeyRuvF88wD/OrGolw/64Q5b23lW9QyTUSjTo9XIMGV9hcDfUyROuf9yMntWV8Hf0uo
rik5bD/37z9OJ+8aDj52YGEHyDuBhV29j1gkASvbg2ddXEYflXlv4xv7Uatx1nuXkoQwnDL/D4Ys
S5PxoSkbAQ8IjcSPvewPW7mZjRrbdHfv2k+i3mH8dGs/H7GIMgef+2MWMNIopFIz6p+Cm3y8C2GZ
U5MF5CyBsRhNSZ29Wmv8KAx6yxpzaDQvGpUbsHPdGrNLQSppjhbXkogQxylP1CkrqeBwa2La54p8
Qf8KisEpjMYZo8copx7I0J9t5YyNfdLQzXXGbZgM7oxuJ/NqYVyEg+MMGj6w6gT0o4YP2PFDTRJr
1iKthhGU2P60apDFJ51pFE70xs5S51OQhKLZMYaffsk/5l9j8s1mQUsopF2A0/KwBJQ6ie+NazXc
xnc5Bh/9Vzd9LElBKM0WjcF9b70pukxZOFsyKmaqW866dLfzsyn/a2InRl3BCsmRWUoRHCaorjK6
K4+T56eDxbM7I0xeyFs2hTlSMtqneVjs7ZTh4cUaZ8kx3sfX6SOsj3BUTWcCWvr1Ktmw0VpgvfDV
RvAEvOIfWmIQzcgG4hxPwc1VhA7Lfj4nDgg2NAla+ICZ3A9/dutTORjLjY4pUKQiFoamgc7ObvgR
fwI0EYq0YXIHiFcooa82BUNyPERDrfOXqw0dp9tyNrmxh6bnSYYQYNMjroQS2vL8ha7b38aBddNM
Xtfmimcv/v8LMIYxqWBQGQ6vMkjBtL+u2LaobjFkcykWKSDfN7wgrE5Tx/H7IZxwkg6b6FCtnsg4
j5qXjr+lUybLodVzON38VjAtIUPBQR6skBDy8+5HMDLCKReH9p+NCIcOm8wPA1go66srYSykZhU4
RRpcxUHCf6MLVgL4UqKKkZ6t+KnTekqQWL63wLhrsIa/fFOzfLqmY/0Zz7q9vy2S3zDMgUkwQI5S
XN1DyvURg+ZCNt6OIJyjvDZrDuNgNL691AR2pUD1a0kP80gknyi2dE2oQcCyFCEkZtmmyeGiO+wp
/BFxX84YmojqMdlu2lwfGiBtR4G73F8R7iSfzrutEg4tETHsHhJAQOAilzRwerzk4pbXRA8ZoPtC
v70T0qgtluOLZykzM4pUY7p4LWvRwYp5Ab/hbXumH5fVpWPzWHZ4kGlt4ROfHJTZIUXX+NES8hBc
PcDCBg9ukMZ+BZLJMIzKsYGVM7GXZsAgC8OE+P+u+lUBUGxv1M+Cf+/ka/WxEZW8vTL8mtwr6F1e
V/Bi4s9MrbsapRrAwCO2tIStQpAeKwCz0UzzGgKkns2lcIU5lgFeu910G0dDuBgCsowkytmysJIo
JWXNERGCgwVX5SESkaysJLo6XOvXa5y3fwnbmxgLztNzT2JCNxPZRapv65XBbIzPW7BY2GVKDFxO
4mFveI+iDg0jJUSOzNOWQU1Aeg7LWl3XFRBuOV8eokCoakzw0AfFWDHFLI+6WeB+sKAg0z+1GPEF
A1z8PbG+cNtVs7MgCYL5mXGgCrJMsyTcWMs2FasM+bS/P27DCwQgF5WjHHMbb4TuHuTX3dcWqXSS
pdW2ifXYDEjwlaKUlCEwMK7y+kMSuyFyrm+aIMrAbhwiaJqIsWGGTUM0zt4I3rEw/uh5GSiwVEKV
CwrvKnniQN/qjAadc3qJ9cnjfsT1JQj0neUbY1coAXFLK9UJdUhSmNWZ6gQHlglDp5+Jb/C9k7ul
VXXW93PpBc6/mPO9OKN8TL4fnyg7G0aLpIkVTMQlPP7jRUT9Y+cBpbOjbc5h+I6hKFxHMvgJ81ow
4wyX8SnhywUrqNvfEwsr2XMHbAeD9IZaNGm5X4O2jkl3/XcTq8DWwBs6sj9U4Pnt3EDl6ZksXfdY
ZHWXAC3efbMV4yGwNJaxb9ArjcC+2l1gx4IAOMINRaNkogf55HnFcLcjWVdP4WFp88h8e8eAFgaO
JrCQS1P7zBbkLk85iAb0cabM+bq0rK3psTatEOnlbWvOpEtO1/JqA84pKvpm7DRH2i0zIiFBluwC
sAsJLwYTJ+O7tDCNU9NUXdDctTqhDXMe5/pFWX/lp29ZDw9nWj4TWW7SyGP2zq3pJEEqAoYHJfi8
S25NEfDLcMD/XdFqWazb8RjvMlPZm+Zh9iKdLrCC0xDm+6xDVD4cNdr++No3e44eM1zRIIZCYl8x
uq/iJJGWrPOdqr1rHMWDDir3wRIAblaG9QMzDDLdCl9QdCSPIrGRacLKTv3bJI0V0srV9mCokKWs
klYnNy/JHzp5YBIShc2zjMKBWzGhdAtz1KcuK3uYqJzqGye9Wnnxj+1QK02wuU3jbddQRO93bR+q
q99RPcz17nBM26JyCXCc+02NUP2iW+xQ6Gd4mVAU22gDXfmMNtCKm/PQMWg/k4tf09/ZkuUCQAu6
EdwV5L2bbQLUTFv3EXZWWkinbL+jjKNyXEN8HrCgY42Qu8UljQkrWzH9wg1Vf+JzuTX6HZfURQnQ
gC5tafw4aiCnbWel6cRgoqBfUY74TU+Ym0hJc97f0Wu83WWMMrTBUBxTaCPbGhz5WjkYpu3qkPlG
jIVXmvGLoT9woleuEqqj7N9CvTCWBIGR5PvF9Swt5Zee+SbILzqoQ6OqmBdwFdLUzcZPzYY3ho87
hPqK7hbs3A9LRnQ5PyHH9wqw7QepyK3+EbsGmvtW6yGFWPFUhQ0DY4SxIZXGA1MYvyAU1WNcOAuK
pjUtsQenkNyky/GZDRjKAtS1k6QG7A1Hsk071vlOVOJ8gE5EOGi7bPqqJsUJW6bn9E7CzJnpehGv
aNy5FRnZU7Fa6mFWvoDnrO2gtj/nY5JvvrJN6pGaDfjbvEGTua+4YBwhP7wf6JaZjTTanWKPcFMR
ZnlvMY6pthCzt8tn3NWowyNt83luH/gdkat1nfXdeOAIEykkPgtX5mLBPVXvwvVE25gXQ0iQP1cV
PDul/Opw2asO4sG3MZYNZOKBodHoyQLR0xRrG4tW9H4vHsDTx1VbvDxQnobF+0SYyjqgzHbJcgvI
BZht4A+v2w8crTm60WvA+P8gucJoIlkcFW3waB24mPngjxDrVVmfxB7LPV7DI6o/TQGHOuHEoN6N
1qeHkT36MlQNjaFPCFM4gpKyYohgISFlhfRFBFLzWvaFUvENBnTiB40FHhEaKSQWKovVCENGSD8y
r2gQmqEQsClArTRuISEFOE0eHLNYK64WzVzt4Cmyf8VCZcJxnifHx14JC9M48tbourE5V+pPXVKH
CP3oUTVYBbzdsn0cZxGx/hkXfODBajaw89WRqPSEUb+FzJOAFDDa+wI5+slw5dytDRwCiC0O4SkO
p49mlncG7dflIKuvI2/mAz/qHzjtlup0ijKyprkJTRFX8Va9nKGIJuCzda3WjyfzPpgauxMW7CpJ
Tf8gRitvYjdFd2DgDDPtIBOcDGhdQYOjcK2fdKthlVlpg2POx/axYYE8XkK2n2jCge0/RLD/fMrh
nHe2gGI5Gc2rg+aFaDGEJWWrWQrGg/R8wF+X5Iv3oqq86s4S4BX36ujLBAEALOf/PCFPHdbJbACH
c6Po7OeI08Vt9q8mbKlYAERjEd/KxHOlk6hCeYHWRoJNV/fJ6mkYESuqTCQIuFW5J6XDkE2yuGKI
EVDcPshu2GKgsD/HIgGdmlU4CC6YB6Of0XzWlJN7FBR80Ty7VAGF8pdmgFRTuJdBcvjxo9BA5VDw
Atlv/FmFA5TJFbzRZLO53NAa3p7+AYCZsmaMSftjgqsmxbleT6sVlvcQp5dgYLtd2eTxeXkyBSXF
bYJ29xYeS+4ENuIL9m5/JeRThyO5EkbjwRQjDnXAKmz1NzeQZs+tfKg7Ozqz9xKmYjPjoFyZ2vad
NDtBLl3opfv7JhHfaBlDri4oGR4EWLNYLAX2YEJaHfbApd0XOgO3bTuxqnNFKyUSVK8mfOJkLLi+
piLK1j3Kc4uP6prfkpAK+MJPWaZxN9YhWmOuPSNYI93rCzk09mvUaK7y0B1MsL5LQ/5dSwc6SCIS
2b4T8U77sqxLyjzapWRTKxc9DgsVOIiU6h+ISZ3jJhReP8Pn1eMhqunz+K/0r4+p5MdmO3e/h779
dCIU0N/UOBo1PCxsg1xt1oB/PhG2QXWYWot1s243agGRS+tXBBJGmkl2VDEjAdGzF/Y59Det0MqX
a15B/ExMRKpddGb4HTyFC/XnX34adPqYV4k140xygJxtVmJt/B1U8E9KuuWFbtjj3PyjYA4kps+P
qLu66gSOmVetWCbKFEizqpI1rISZ2rrhAuc/6nHuj+Xw9No65YqxRRUT9qsx9VYws9hLvNXLjhvE
YfzvAqO/6Dda9ugBPZYnnYapnglK8cRs31R2l3xi0RNhxRbQjBQ0gSCcNy+EMIAICQXx2xL3ddxD
nk/FiW6+wxkaQB3NJu9LOVf0ZvVPW2Ymvt/yFcri32asVb+33kB27J44nfIbQSVhRSUwuo9LwyLj
/edoAn91L7E380WAN/jXgzKvYiQ/osnBzYxAIaRkuIavcsBUS5Sl/5aOKHFad2oPrYCKRlJHJAGm
VjNEWQEGsXyk8SKZf0xqqWPzZa/w5Yi0OFpRRy5kYAdjac+U/c8cJGirtSbOg9QIEFTHGtT1o51U
zuAomsPBaK827KZOjuOtgSe9KrPslcGnlzUY8O1LtZzJXRLXo3liZMZFoD+SJO7pewE4md0V8ht3
1xuWSVAW/Jw9IP8vVc1NxeOqmimBPCsTY5TL3Zc/Z9Hsku7nGfuiQJiZuLFnkRbhPB3/6btpYAU9
oJ0JaR/ax460VFeWS6xTtz02Rryc/2IEK3/taBOkkm+ya8UQT+clyXkl+vmRvK59J0Vu74XNtTOz
3r+crMPYvahGnb1RKArvWdn7AYhfEgyExR74cRd+t0kW8W2WCeuO6YkBZlQbCyaKGNlJEad9GvKe
GC+vOl9Sw3jj0WSkGM9cpstkzsIJgzSeT1RMv7M/y/srbFvCAmGhtQOFldwgzCj+Fjfcrx9y8tX/
VCgPbH+LJ6n1+3+kKv3wCNvQ8Ok8KTEO1iXTXco+NeDlYCksGMPAtOj/1ozPq+UqZDfqyrdwK3wt
g3MMTqZFANlaRQiMIg/BtckJY00QhfD+WuDlukVFCkkYvvPjOYuIghV48CHEgcJ3u5Ek4GPcxZJG
uRFw/xmu9WBl/m050x56xFHw36aNcKrVgfm7k8hFfMn3r0u/kzpZ+sB10qB/L0SyMksGK+sAIuY5
l/nb/DS3P08akeDnGpwfvtUzCr3cFUW7d0Y7cWJ1v6E02aX71RukhDFQL/bFEmC1AViXAltbXbWd
+kIRBypAwCjp1idrQx4HbPnWwkwnhNfs+s7M0dm6AKCMvrdxkP6itl/9DhDoWB5npeo4nj/MsVEy
Me8MxL+f/pZneU5icB0rzuFfSEmHS9bMJkFzYpAgkmTBYrph3zIw91tlVAXWBPuM2zpwxBEW6bti
9Lr/j/Hc8kCcE/qMDkC3PfEMnvLMQhX+OxVHUGyP+XsESE9ufBsNxmgzYXC5oiwiuG1NZH/oCi22
x5aE0Lyk8ck5kofhnt/oQp4gLhh2esj9QhFZFEKArg3JEl4MfI8kVW1aPXkYlumA6cAsFowjXVTk
dkW1+9cYgcq3FySu0vjH/XkKf5cRvp4M1O93Ms72/hS/GeFRD4su0DmDVm0DXNcEI7EIEpBqvn9+
bkP8nWBHoHSyIOTu/vF5j3HYaT5JTt7CJsFy1ol4Ye6J67cub+K0aTTuv450nVomnJW9NfWsGG6K
dXuLXmePzFZ4u0ATev66BXLNI7108M/AH+XO339ElUwllVtwhlkkTH5nl6flTFB7nihjmm36xOBM
TEJr2LsJNHMQROTMRESNLDHyBx8N0De+WEGADoMGLDKG4cT4KsKPNJ6e8yh86KNeyDgj76QByGyT
kNUfRSA1JUmbuYrBz0ZwhHiSSyuMOtgIiwyor7mk5H/J/e4JUYMyNWMnfr0kyNwkHDQbjmNfs/oK
GGDeV8mTNmgrOYGV37D6PKEiM75WA1G2SEti7vooAuVVzEKkBlmrCuQGNHmZJsJqZjqkba9t8z3y
jmAb2itw9oQc/3QYjTnObRMpjKuBG+7+pJIcXuC0+52gSV1o5qwR/+g+KrKnuXQewUmYNutsCcgu
ZAXlcEHPxoUzuZ6bcMCupihOju62XzN89ZltxtmpZ5cnEIt06p6mKpAIU4NHCllMsMXYc+1C5QLy
UW4T6gQpWoVT0CXqf4EKgoa5DceN/DMa2x9wqiTxhyVgv6y8KdIERzkERtnUqe174RQOOL9Hottl
17igC6srI3y//vVySd2amhleC7i2CdUaUmLaGmvo3NPKnuDwwPzi2dF3OryKqGu6NAZNV2uHKRNJ
afcH28o58r2XhjcGX3EQpOwIDl5FcEKG2qN4OAE0cqKFd7VOpKzH4rDyk3K1SUpHngGi3kMWyXRZ
y6mdiio204lNdvAcTXGKCf4g5KZAMcmBg1+r6ij/gjkqYUnlIVXJmErPRBdPX+U20XR+Cr2Z+e2E
oNf4xpyabcj4L95Nf3pdofXlEhuc3EDhv1MJpQ5gnzv/zKsYFJSWGEhUoVek7gAdOB10/TbgSH97
wMEmcx70y/G2MeFXID5491B5Qz38FByWWMMRE4eTBy6x5Et9NudcR6kjYIjUI0lSj3uBnb/w37kK
V49KpE0BJAuKOmlp4Y4JJueUjZAhsf7SB4qTeUKt6rml17l/3PTzUEYRR2U2CJIxio5H3tEVulbP
giV3Hh1cDyfv/mwbqzabhgAqumcqUlQZqfszC4GrrJHL813qeF+92aU7V2Q+J1jc8cBaEda5lPBg
a6RGObomu4vIbqReFSJgnmpuXr/XW6Mqlciu7Bmog88z789ANfMUSBTFVG+KN509V6ws8ywfisIX
X/nTxNGr9XG87FZbNfFe/tjLxFYoeg+NuCRWnTbv4aebzE9KNFWymfM4PtM84jw3SHqveTl2JsAj
ZHp2yMoOnbrWqCvTPFcdBou84LwXQsffchQ+08UL/Xv1p2tvzKC071kp1ggIHffP25173HX86L7r
l0z48teeuR5WZ7mIDr1zRnzg3lfCGYzVu2dWaV1r2NuGE4iUeUNX6o8ZEVP/KrIggUCcYScVLuBT
W2H1YtddH7SmFPLnUP/ChS0x0oEgfoKMeiR8BzFM1DlSrv0DDuNDJysDXXe1bhTY8Wm5YidvCHOB
+Y6YLmMFAJySagelvKU3kpOE5RosiFXWLSymGxdeDQByRMdr5WWv9yb+mXVCDXVxiq4cvSgjwdmZ
WBzmvOG7GfhhonDcSVpiwTa4L35yald4GRAn37HpC/bkVuhGHXIHGq7W7IMFH+Xg21YJgRCgFi5W
AlhtQQxToEkCmHDUkZcgcgArqgQIYQClzJwxGz9O92VQ0oYLv7vlonV2eOfyceyCGDsZwYDvFXa6
Z2FSnEYyA0/pzF+gwhswUCZKeVDGMVwrXYOM7l+vb4Ijs+gC5epCS/FXvQ9DIMcvU1fZu74yxdiN
iEZeFiOSsuYdyASeJZ3nOk9m5oJQ3XBrgM2IHoil3uZfkRTL63J51qbOVUMtgH/Q6ZJzXJZr4314
rEwZF8JjbAfWC1rKaGCG/DXnNsULWJTWhrp+lGmksCOKwnQ8z28kTZFza1KPitK0Bo2sTQ3lVlEO
47+euR0uYEkz5Vf53aWOsmqtRiXT398G8osLVE4i2+27qd+FEaOUnQ1YIoQUwDCN8XhjO82KterV
iZ7KVPC8MBJCRhHqczF4LqqBft1jcABxsXLER0hxoY8oQPjR0vUNljCdjHRDk/89PAFLSIK1b8XJ
vVgcSjILnp+Mm2VD2hGck6x2pxurMiqf3Nm8oZLemvzCOAXZIqcCPBzOcQUGuo69rsCPOX+0G0r2
fp2eMl31NdOichd0iHyd855qEyavEWLx6h/omwPaHylAr4ra+6nK7QDy1mrzlNvevz2kUeSjYxVD
cJtiCkqYEAScBAsHiNk2yT1wOyjEoTr0tfY4Oe0T6KB5LMtgfeJvypPNRYOHbDXWSE8DdHJ+J/gf
8v1mwrCVWeQYEhYENGAK2xI+Nm5lfQTaL/cqOMYT+ivpPOWh0A0j3NveQWMxvWPo/oD5jlW2njgY
fEbwICsrbTpYlEvQHWAVO7M511Dql+b21gp2x1pL519cvbrfptRlfvsq4ibz6kh8qlN2+pyvAvAW
OqHWActw2yxpTy2aYjHgEHHTxSgkhFzf5HIiqbSFSrWL2IGzjtgAwvuuJbixUMSCese5EkTGaOiU
ekrgvVR6pvwz+SPYtQ+iWf3uZAJslR3HX5x9wXHIogEfqVKC5xyRYh0g6A5/WHo2UfWK/NWaY7hN
KBNDGfFgO4vbYis+rWNg4PYZdFHG0ERLdXIC0ARvFddVbmoNgfx/UIUOgJwDblQhcdq5xJlNjKgv
lFwfvDKvZld8DmytcYvxS0e7ajkKMj18JaDP20OZmpD3tTlewualfTqyNuLODl7YmS2Aaoe2I5XW
C0mxRC4o2Unlm5FVIK2YR3rw3XVB87yG816AU0LtBglY9+guskqpS2M875yW0qWYPfciy+FkTgsM
zln6jSPiv9rXzCbjWu4TdgbLonMF1z88EuuHlWI9+7wJgiPTMzxYtHGSkdbU/JlJwDUW21328E5e
N99QW6doQ44i5X4qUU5PrA9ODcZLs2PQ5Laf0nF6v8SSn5ae82oyS52w31CEsanM2e29Q0vOKM/6
Vwl08ZGnpSWE7k1RVJdTi5fJFhk3ntbW/sWACUD1CxVLY6QXtl2UdSrqbD2QEmq6QkFCkxCb4dcB
vpdlIlBmCh9VWOG5F7cs8k29D24NOQyQ9jtX6Jv3rUUF9EyrqmiEvXDyNRF5Xtwng6ROUutU6XUH
yor3IA2D5nqeFfCaARf5g0w1qYTWhF8pzWkR08B0DQYmxAw2j6xrrD5BvjYW6q9bXhnrvGeLxn6V
DPId98OfVEvX50BYfxZ7EgPOkVX9VR5NQ+7DHQppBrY2KlN658xN/kYbcoZ+hBA7HKYumMbCx2Jo
ZtOhSWAcXyoSVmpcGEg2pzdZHhT3755e/wdmcTMrTz/rILaxWCIZnDxdvnmrKxeWuVguqUEjpkcD
VafzSRiAyjn7j1Yv4PDO6ysK4Dm9HF1fOEpjrdTQe5/q3geCUKFUFUfXDLHP7N7C7asMmWn9sh9+
vICAGDa+CaKqg+/WAoxgkxtp4/FP86PQzzgA3wOMGaXHPn3UZRnzxXnP0nQwbqpgVJd6dgOF3Dvm
59vpw7YKzHj2oEU3xE6NHyZnGrpijdQravM5BepA8/MazZ+RNlt/6Fiq55jGUAXmXDELlPfgJ+8m
PUHkyEYOg6ELrTNwqC9FgZd0WbP1ATEb6Mx1Er7Ht8wwoXL4y8+r3yEowPw0MZ885JGP3KBN9WxK
4eLxl+5SlJBUqOJClKmY2dBcvg2Vce7tQ5AKc6BoyAgoo5fjTZYWMcgYGPbfaUvFjIwV4r32lTzA
TX8OPwo4u9NPD1QWz8qn+5nOEjls3eWgkTScwB4kLsMaOV/HCK0cHjfHoNQOQTplmIS0euD/Jy99
fG6mKHpqMzN1XUy3Z0BUxGl7bJt4Rbv0+7GfoZkosX4Ak/Te8F52AKqg0lcbZidXtJtc4BxCSJ24
m4UfgaTv9PH099fKzYAncAJYjXL8h2VQAwO+7QdHxDctmJn6fvWjNrq6OayAOe9UcgMXKDg1Mdsl
nYt48oKdaER5ZF4kqoxv9OBylVuN9By6LVGHG8jqXW2GROtKFwClOk1r4v9sUMjwXIuKbpPcmgMI
BsEfeMYqyedJKHDqfdUidfpEpPdleL5Jeb0wWKttxbOPm2jv0c3RLp1hu4ZURw1DAkGtKh7rql2o
AIAExU7XKlV4flaKI6g8o/6rT0fVk5eHHLNmmeWZt+EPVF5BUGT2hy7AupzW01kQYidYLdx1QApD
fdwsWD8Z+uj7oOYAGFX+y5aGFIS/U+nVSElVMWX95DkTpUdPL+O4LmEIjiVoYDT50d2hkeYmlpOA
oQE8l7rC7BPNMaNthV+fMRaAb3NZ/Qrvmz94Mq9Y6Gl/mN4pJuN7kRH9dEolS6x1F4V3JnO5rXDX
5E+Hfo4UsqDdwJAt/rqaXhsNIYUeJJpH29ewAZSTU7r+TIDWNSC/mUt5Y002q1NTJRryWXyuXZvP
UwgWgw6J+Iuy+dcLrrylZg/4ousB8cEvqTzOtFGB0127V4eaJTu9PLeaxdAKHIuR0YhI131+1++r
okCaor1nN4Jqje0QZOsX6v2qij6O14i9UEhE4KU2n7ljK+KW2+sVKQVdjhPakgIS20fdujm9XDUY
koci4pnFFwzXegZPsHYGNV3HmS3K/gHksI9A31r5YtfBQoRwc9qmjRNaN8ELhJmfrtQMJPGxeFiH
COeQG7FafdGNooZwPAldPuwxhX4A68Pq2SCE/tIUjDRJ/dxFPx9WNCRmxD2jcLeJ9H2J3rtvPwd8
5LSsTXQV6YfY6rtc6VeiDLKt8BlX5HiJsMqWOscilB1LJw/K2gZx1ykoXHO2ybUYfXo+LmG2D+CC
HEdPE5/fLdp4B2B+Sm+h8gMC3tsQjhVPjbvP3ApxWkjuSAW2Jh7N1oT1LwC3Q6Fq8EWEXVbv6VyR
FMtX3yXrUj+4oyHaRghOM2a2VIqN4XiCVZJwYbt3iI5lsurUQisDUoMHR0/EG0PJVf3ZFPgwzYrz
v3Z8JH7PfaJ5FUTUvTh1lJxmB/788Hjza9kfWM32OoDtuPJFheYigik3tqp2RLABBV0uAzQNMCu1
JobwJCoRE7dST66c5BjR7+kbEC9I7U37IRJPCgoZOxH/Wyb7R7GWe01DKbMqdKgreQ61NVENLFTg
D7Mr9FR6HzpKC/1Y0bhjSRGpJc87YzrSN/FwEi6zyDj0bT3NzRU1IojZ9iXrExoQZ9WoICVEOsmK
E4xbGnSo5IW33gVqcrBYagDPXSzIzqSDGHvxlvzj5bOLIcjORvQwgx0lk8OPi7D9HmzIElhATXbw
YOxLdMn6ALmzi8r8m1dNHJ4TDzEXY/cYQvOl1daiXjzSwNocHAo+yNlmbi+dmxKNaxvu92yCgxV6
r+bDBmnX26fvaQlLq+6bpQxdCsV/qr5E/A757VofYU5ILZ2H4OJzV5RI4HGHrS8ewK/BwOqyWrHP
PcSb/z9f001qNMF6jhdXISIGDtjroCtGwCLmZJnty8gjfAiZ2Egj210VT6K1ESvS7B+dfuRXZMrI
gt3Eebm+pwF8wXGSePBr8a2iIJH8z2RGJp78wCtPGBWgYvSrIgtL/YnLXP2yrYRndomJOQDXqRJ0
8HqaOqjjrAGQGDk133i3NUQCyQStgHNxCdqW6xVx1d3P1DEoDWPgO7pQ+X0MsCWszCwO2Es3mvgF
nhOkc+aHuxdERBevigmMrcPy8kYjknELlfZ/74GmGYpHRLPVvhLhyrt+9F0kwWwOXjvPHFPmruoa
RyaECIdMEpCYBnShcmCJsGALs2MT3z/DH9pzNHw1QSH3P+6MD+1fE0K+2Kf7V7DVwmfjjyJaEur4
hB6YvYJ0bxuU0CZ2Lsi6Odu6jkkPJm+U02KtnQP5K35w1x2fd9b4gb0VGaX5uPWwINm/x7l/O8D/
TGoWXh6jDc8MkAmyTTom1g/Gsy3N1CT8r6SkVvo3RVTbAd2tJzsIX+qTO1cuONRiv+s5M6iCI2B9
7CvD8dkMX3uGb2e0ejys1vd/hoVpw10fhAIZUyj4UhutIsSHSympBPcjqdTJOPEm5NIKNK2NFLU9
1vTxRv5zZUY+2YiI+ddLM/12p0ls9m6nu3mbhgOgcdQU+RhZmM8f61TTiHLmnHKAXpnzvR+/YoCu
kPwMYqc2XvWIjbNqYTysxs/RtGFwhzNSo6NkShgOO8uVtXeEFaG+pJqGkgplYh069APWr3u/ABO2
7NgSpe3Ysv1De8z/Np77CP3rwg/i4UUSGhtOVJMfVD1vwwxDQSYbh1VFvXD14m5IB1ur6f+hRTMd
GAKEWhw5aibMtwATTOVKB/o54jNKyEso9IDaCovvcYi5yUyVQxvehqlJ9fdwKx65FV+0K69dlBHF
6viEsX9lL9gyjwpaOHPvIwltiOuh/9yqpvckPaaUk0JONLT002yKjQ4MJqdzl672Bmn9Gb2DJrbd
+YDtrTNNIr94e3YolLZlciw6Y1GU7MMZALaFW483RldocCDuPnNgD/GBghwWVfWMTAEMJJ7GDxbT
xuU1UjnvDakWhp//bdzxN52Uemk9CmqfFYP2YXkMzLhx/rECoyVKul9h0VFyJ1IZTZOEihZmZ+ln
xwAWD91HujA1Dc2ckbHanmXRTYcypz2QPzAdpD6N+olrgbpg1RVBaTr05BJ+0a3A53noio2ZtHF/
GV0+f82ZF2HAqvgugF/rhKTANpDMgatPWZ4eeB+yNLOjaDF4byYMneyFnBdnCS0MHV14ELj5twQj
qo3YLZGC9vbSCbEcUHX8TTTD/Ek/UYLjSbzqEaXulArvaW/FWqmsGxXEsvHmKxZIquLYmqYtGuvp
81XWad2Y8dixOY4+mD5j2j6/pBfFDBB338jJ5SQOIrs3EokpTpV7UIfm355CZpzDPb0G4/bxu6FQ
tedVGsh3rGe5hYgzTKePB463ubSjGqRdQbfCBGx4Pmfm5/E4NI/tzB1OvqFpqwv7FJw9JkIwcoYF
nr8RYxP//RXCeou9X6c10bslYaGt4fAdrmbNWCPQT5SIQ2CAUdG3ZMptGu3onpGIEbBQss0weso+
ofJ++E44m2LQnUUWftvnMyUpoIQJNyI1kQ4qi/G6DYCwVpyht2uPX+TNYzNydQ2ebzmxMGQEPjGk
v55tjYhNHYmKBENvoOwCGGAZp1OhY7Mn+SyjHfhz/gTncZ7Rcvz3NJbmX8GDTf5q8UUkFwNEtIk0
HTIRjp7ovVYJ9YA9/Xi8JMLvfg0csLYPHzkZksPyf5vmSo+J3GzsM2EfKMXufExKwiUxkUaawmcg
0N9YnRyL6fX7gDDPusf8vK0F0WBGoaJ2KISZMx6YVPbYyTZyB2chXsX8VKCVMW/NUoDju7ANN4NZ
euCPkyk4P2iGfPZYcleB2W2HmsvtNz14MJmyV1+0XLODcAxHuGNzTwWehbyNowa51WY2+57WfRgl
h6dCjmNgfTEdZ4djqDCIhw2IaOCanZkhUIl3W/zKaW4CAY2HvIUONF0uEA8LoKRYhSUUWc51S8Jd
2/SPpwlf6BS6+MWPJmjc8n3Fn/0SbWmlanYZAkTkyw/f2Lgf4ai4MArZf0KWqztT/Lwjl7MiPqx2
llx4j12+sqxKtYZjkt74hznF9h+ufgokU7X18Vh48oHI7Kyw+hZuTOM/5cDjOXe4vyBXdQ/WJpFd
Tt1uRl6n0hsVdjKPkijYV2c8oSyIXtAbLdeqkVvZ0jyxTUsead9xlTGagB1s9TUBXTvmB6EXPJgG
3Rr874RY0wXaMdW666ywsLiV6V+Wh/Zxf+2olW4DroErXxF9bGIuagX2iHDY5DLi081/zRtScbEK
x0oKqk6rt1s6h8lcg6GHHMvQXPLmVwf+6qGj8CFhlDZaokv7ZsylW1+r81R2j6AZmw6FUEiZWV6i
eykk+V9Ips+boqRDBcO1V/8ta1Vo8Q0ZgSaQQuR8zrnuCXwkV0vO2OT1IO3ftDdisCPRoEhiedpt
8mNR8fInN+dDfZWRIHz4PLALReAN9/h6XffVn086fbUak5d1R2945cbOm8DNubDbJaHs6l9RAL3Q
6ZFbQX6nRcjjfpSBncNLV87QcqapNiiUowOI7BeJI5Avx8j+pZ0wqx+CD5pp3vF1jx5X3GhobfsD
TqghygLWZmkZjgoXv8Z+swIdlaP9Th+rF+qxJ8c94efgisAz5pSUTYPkNgAynRDnwq+kg99/LuCL
fKSXRnnfgwqKegSAOmiNojhDPyi+61n2MRt1qry+9tRg58kLX9h05owkDUdWsWikC0/coFthEf8W
TwQYVa7wfn3TRhkGNSJTJVqjtLEipckNYzSGM2p7P7x7Y5fvm+DVc0t7qVvE7GqLFTktjYEXu0GV
UEJx/IwCwSv1tneSYhCRrQCaQU/xyi6r//r5Iak5ASQKuayag/8NHKn4YBeeVYQbep5il4VlUAM9
VN5xFb3E8WTe6GrHOBfvao20D+3nUmNCi3P6EYyQjMFKFyWnq+44RuU7veClMSqDbgfnCW7m2QTT
BEZAqO9Qg+XLlbTy1VXza3hRLyXHzkmcUl/GyacXuFin7srnkabDBoN3kOw54q2XJyDY8xtSN/0c
nrdbjy0vHaAryzKCC5JtowuycmPqozUpH5EZ9meR7sEr6io8mowl67PYj6zhqKXCyLqy/I0ScPj7
Lg55FtXOeUQrZ+gr6qLM7T+5ZEX5teVPh62JiqBzGZZugWxdRTUjb9LVvF7EL7Yr+oh0evZu2adi
DFtKNVU75h9JPDRuvpT5W71FdtYJywMwlHxtS7ysro3KaW+WXHcIulCZnbCpOqgex2tLQ9xxvqSQ
BiGO4VPgBML5/ME6U2d9F6m2MayUntBdU7VY0oM+o0lN2NP5S73lHh/OdmMYPxEfDZzcSTs2EOkI
UfaTWoOQvmKxVi/KWKM/UoLqAC8WYH/ZNIMu58iTOSPT1bMVLnpuPiIbyrgZxH/0A8PY+DBPilWN
yP8/y4Q27CuLzx1Z2NHW5Yrhs6wUkxSa6kmxgT31O3+GhEEBqgcDX2b8vLjr9Q6bZie5LlJEDrov
dwwVO1dc1zfIKGOPXCQgzikqk1De5H/Spqyq9216ohATG2BtvoAfI5XL5cbCDKlQhb30+EhBlcTS
V3x1FtP/bYmy6jQc60ghNhz7pv0rcIyUtVFXdRO0JlBOgM5GnJ48vxaAVCC8bZYxCBitvfv1E/IN
b4XRUqVW+fcdzZ1VvHBtvxwss/0wxcn640IGPJJ207SLH9hBZ4SuToXTS7mNkDmVoR0ARj2qCeWD
rkQL2aI4OUjdS4uewF5IieDIhzexEbp+ox9KxtGvszwLThglqJe9a8kW0GkEF88utE1YY3iExqaP
9fj9Jnzp4BKF1Sl0T4G3X4UlMWTDAR03nTVJ72Zu6N+mAiJR1yAjIERFn7QgGstmJNXN2N4NHPoH
IEHbK/Gq/yafeVZC6SkhrGUX/6WWH9LgJZ9zihi729+9VvAOv3DvzrQU/BHb0HIaJzdp7KsT4PZr
jPdXrtnjMw/DpzpkLmha9VXC2+PpLQj3A6OmL5ik3VNtaXNM+OFe+PGKuS9CyJnNWsvTtpTEgFje
79C2JKU+mzg5Xjn0ujsenNvX0zwP8b1B31nZ4N4RGKpkvDdYV9m1Z17YTjKC44qzp+OlTOHN4Oir
OTdIZU8PrfnGsZxRycXXop8MWGIf719pifi+3riCV2sCYIxDES4hzNDz4qqRO3xZnWEUwNOCGRZH
giLxHF9/0qgvrwMwBitVW/ed93PM725ISnyWVMUR1MSztHBL+k8OBKsw/sQ6riyVjgjEgpt5IGUg
e4l/d9+GZdPyvsdzC/qiWG7g/4ka37zsKptmb4psWin5gP+jUk7q6k0GxmE9SwpABo0TfA23USfp
22TbWXKI2nGIwYucHRAsAsFEEEaeflO+S3bzq5ilV3mdOJtPlzlluJSWYMme2/1IhBIFDdyZLIHN
gZX2NadzrMavqSMHrHLAqPjX7PzZqKl3P3rqlX8n50daLhU35zp3Uojj9e6UiVheNRwkPJGqiqAM
bMk/L4lnaeYPLJ8ov+XzN8htButhfwXQJL3+Uaw89ycJg6rIw2AoAImqg0sKdeLfFho4vyPNEb4G
3asJeudDJZ8k6z2cE8z4xfxuWYRtNPlyUN0n8awf/iEmjlwmofhmxfaJFGNj6YTrgA0BrembZ+qG
hD0U84VSZitH+3NYYgst2K3mZwpgnAzjY1xsW0JJT6H/4m+QgRNvQnPOfOgo+3wyhmpm0oONY2T0
zzKsQlnSGhqbEkzcwdEdwFK1K/tfyJBVfKhzVVH8HYHEt9cpoWCKdcRrLn/PyNpHdy88RBArlQY2
qkWk28OUxqmydScD/Y2nhGTKnJQp7JSA4W/HdYGYn0gFUJ9z4fAq1/25OBsefUiAb5sSM0goPyvW
vqEC8DYnWNSIX7OrIcXg4+tmwQVKYHxKp+1wEeIm5o95IYNf04py5TWAX2poWrc1fhmlrmJxJmvB
wCAp/o46LoouX5BtstgOiAiMhFhQmJFQZxz0RuFilGfJTf5fRXAOD/Abfa3TtCAYK++wegWTH5kJ
02ya8/qZuqwSoFR/rFHOBh/EZHnwOfaN9pYPR/Dox6uWOqG+5Vp3iai53uSj8kI27T8werXQFD/t
+7ykYVfHnGDwGrFrEWGXqSb9e+3XMhaXWevK2hI+uKDlJoiYNUq1ysDEba3xD1ddIZbl5hkvp2Ut
h0cbcRIGAXe9mENUUCS3LYh3u+xvMBpQB8/ULB6FkZQhfVSMLWKkuxETF8FVUdR3cwME/IEDQ7b/
oKIkUgjPx0z985CK24zn3nfj/Va2ZHG2NtsJQc6H+Czv5UIrnrM1M1dZWs1bdomS+x6P1OZNzu1B
8jmK8MwZAnfsKdw3ddMUNRVv/yi1ohceXw8g91aBf2pmNnWSd0++tEgMCcVmbbde6Fre0jX6mEjc
zaSzDQiSRM5GY26zooNUNUBpa5yyHmOFOqilCz+TRRWkZ0EoeB6XJkiz45ss+ybAZ5fBkp9RNlBw
KvaX0Xl/zi2UWXECpk4hThVPq7wRCn/gWgVHpATNmi/vhxGQnFcaC3ep9K8OCdKSlZu34aQ1AoYT
vI5wFChTHDyAdiMOQBWTjip9Vfe5J9T9wwlclYpz0BNTSKFHDrNjcx1N9A0EKuws/I+8+zgezAfu
LurUS0j4/8RmH8ciADi3TKZ0nknjeflMBE85UoNR211Y0GcBgUsps+rho0MA99kUIHbcbG7NJf4P
zh2oUkdKnQORJrz9OO3+CebxPzz3pyh39EQmIngoVf6Wt7aRxmNu30Jp7OvHlzwD2Y6qqK++N2+z
QtHbfHhKl136GnQqMHyrdGr0SMPK8msJnOaHunB8pgpzNbLxx4slb1zhrV2IyUXZlxgKMKGxm7cW
U4VIofgBC2EfE1gB/BiGOt37ZLymEIQ0CfW0DI3Mw/zPDvp9VdRQs4QFm/H3Tspz5Hk2d+YEMww4
iDQDI+SE5rlbBEhgAkEUa8bHSWB/bE0Eheh2gaeD8zWLUNNAekDBkA15dcSXUHZAo5MSGqBuwte2
ITsPgts63NvVNeegQ6+CYhVDtdXWy7bvpi3ep4jwEikf4Bsso3zQsImKWCjfMTJeUJWViP2DsR6q
w0/LZaTPos6uANnSjSuHOhz554zeybrB/PGngjobK/hruv9Cxj7eshsWAmww2izBV8nA+Uu1nDpj
4Chd7npiYyYspE6KpNrM+n9wnm20v2q+deMgjUSzzm4sKv4etnaO9WuNo/qfnZcobz+b7YjMxOy8
IfFWbPEsz7BkOtI3NVUa5qfZ9FUJB/t4R8u9nNt411vvlnOKOmZ72sZO+9tx1bNGMyXTQpZiw/Xq
cnLopCuNHivswZm5VQPNXdRV8ciCN3mwQlDLhmM5cUaGi6u8LNuk2GKG5H6XDgCiIhr56IYbcT3d
6IfdzNsypx2SVNLpWinVdxAqj16o6KA6dglMaNFa7WLHY0U7HAa0sn2SdDwNylPFaXaHhKvxlIpv
S2K2GbL571dnLv4ofufMlw+QlBLWSEga3QyKS0yjLsPPIXqoRVRlhj8W7OoVtQbCwuGVg6v0n3O9
MWnpeo/I2z0Pd+2ajQdPcBPX5RxiiEs9iwqJkD7lrGS9IAlPd1aLZUGO/i28yPTdN+V4Pi4qk0oJ
DRv77FymsK/EFG7aBXRGAUu76znwha3/kmMXoYTXVD+gBP6WPrHj8CySjg/wO0Ao37kaRNNEsNjK
mVJJleBg62kJ9KFPq/ZD1oPj0PLIVdllh5hkqH+mfghpE7Zao6mVzlesPjIGrqbf0tc2bU8HZNBG
u2JoPNSec0wFKcliVyZ0zTtKqnFUlGwxJ7ZvmXw8L9U0/1bswVG9DLwdaKYGGk7bzH6CHL1jrhc6
JC9u1UDgtz/lkA25t54oqYCJ7aMy1Nt2TRPxSAldBgltsnSsq6QSaTykS7s2j5fqRg+5qd8RbU8x
RX6miRcLKq2ekEaxnpu4l5HGMZ0gP0yT1YnJCj3QnWEmGbVFGQM7i4M9a2fnUZysOxhQQLSwPQds
sU8pcmLHL/CGH5EjiwqX2fkJR9nyfVgVojOzrmU/o/bwJ7k6qJWxZAJRAVCxlbNr3QDp4y91VWAx
wLCOiPpTdOy8+DXKszL98L5m2BQyB3VG8R8J704p9pdTgVueU/mRYK9BdlaTNyVp+sQ5t5wGvXSa
raHP+F+D8n8nHPKG9OvqJVOhbQC4IjiOaWij3zf8KgEjvKYD9+xt9qGKdR6QJ/HHbzxVN5Ma+6wJ
HER2AxkB4iXFPHKDWSm5YqEfmvSuMKs2JN1xfP+3YKz4DFoJCBySxy34Tbu26Zq/TjHrBPBgMsep
dOTtz8gwRs2tg9O+dw/VtXeEcYC4OqxbzEUO/itsBQInBuUKAgXoIUpGTCB4LPFFB74NGtnUvVCT
74TswVo4gJvtnLUo/yqRhn6jtzfuSpDfNhmQxrVIsvWSWLBlzyi2FR41hXYO+mSSJx257o8Yft82
GyuegBu2cttuLKwanqd763O1Qzlrgne6yz5dVQ5pTMifKe3RLpZj11KU6h3uKdVjYJtXAURODKbE
uXFDg7hg9XqYsaOrMme1sSjWVbJl2ZkXXCYezsZcddLhp8PWLRW8RIzUbE/fsB+oo29REjmPsn7T
ZHSQeoPdmHxJb3U+whRpL5YVkppwYSTbT4qoSKp2kRVrFqb5QfaDCimmRTgaUKyO6QbhLafIt5yf
fRSefXbn5FXPZWt15Vl+/dT6Sl9yQ1ZbLULkzkmFV53ZdM5JLqjx4bFfrI5j1Xlg7QYirwlhyIu1
7+JYZ0yZQwS3QrKVKyMkPp9iJZt6I078m8ui+7QpvtPZNyrjf0s0+zZnY0ybTvpGaLa5Mu6VeLOF
tyttMoHgSuSpjFY3D7Dke0U9y3UwPtWbDx8HwXCr22QK2IkFneSrmWmr68Zl0rgMB19lAjiB2ogq
oesbtGwO+t+JRQ0i+kk7qBFuF2FvF3ts7yeGB+rDQPFIrtdDD5YI3OS8PDOWdXKxVcWTV4BMdA/8
JBHmRQU5rAJ6zaVp/pwyKKEZvA62Y9jDZQG/0R00OOnoq/XsC/JQ/1sm+x0/+XzPc+JkKKKqx/vu
zIiEbC1Wa5j4E1iJHkSgdnJ8Phw9QFqbb1APjWo1osksWhNZPygAzgwbALSlAJaSKrTSBWtH6aSu
h6HGbCkrlMByjYawdOq4N4VGzEN6DXdhiA8HOHOzdPPsjErpkeZ/we261GRNaOcpfTDCycPWW1ba
65/OJf4PWz788x2qM6De36ixjsrGCR6nt6FcpzKJ2KaX9mDxdLKOH0XGK2MSBIO85qEz+XDV7s28
9SoLnpukkAXQKbjGix5f7sEF+gzW1MTDof6aa18D+s8EO5SETwEE8xnbWWuBUzCbBkBOJVLxUt7g
7TJauYqSMxWHMjRhbEiWm0qxcnyWtb02nmNSs5EpeQ6HJ2w7Y7OffuM+bY3INusB80ioPTeJ49FC
KEqGmR+4QFHetkLPV0Rw3n7ocK/Qfkn/Z4SOrbGkrAmRXfG+FDbx2dsHzAG6L2X3SmwCUrO79P41
kdB6dQXc5kru67vI1Vd5z5lAIazctzDhpq+SbPMJyn/eYI2o1vif3LmWj0IHO6+srpRN9NXRiq0O
GwKkiGkjYbpak7NBT+iATFBv8BHUdBXQF9x25Cfu3RNcEgpApPwbkC/CO9s5kSx6HXQfU3s51Q24
jBhm+kGwctaWsU8FZGxG1m/ILID1bH6u0cCtK0tg2c49+zthyrpEHHWjViKETHjMwt/TXKY/H4fY
+gK46g8Vcwjn5gcl9pzh5YORArAxU6Wa6IFpXIXVdY5iSlsZPD2RdTh7uuxpjjbpXr4Wpk+aPdKd
49YxCLgnD1aGfsqTYKawxLPKJAyoIty5E0Al+e2ho5/wg5TlA5TD12H3PdU+yKBqTwOg7eLX0y2K
L2HaXHTCbzTA9rWcbP+lAAq9UO6KrBGVxQoXsucwnk6DaQf4p3NSeaiZBuvdjag38Jb/d7WcdctL
i+QbMK3boqkTRMK9I0YkEc/UkpmqidVjKQLNzjoTYkqP/tlKE1DJ/R9chknRm+v46PPNTJkCsIuP
G+jrHbWMOsLBUZWU9aOzaIoM4drKv2Yq4nKQf02qJ6SA/BYdJ+SV55OVkEraadSx4wF3k4hGx+Ho
ZiNiiaiqVaM8hzuSpe79kzTZqB2Cslw25+Hi99QNlITzWn8gyczXJZtD4F2FmOp7bHyp4zXjg0nB
qS7qfvNJqK9Alw3tM3XtDHZuHOg2C2xS6dA7jXS3CrB89UFcYyv9rEprJ9BwKaz4JaUQmbHHYmw7
/HuEu2Ipfh/iEIopcntqP8I3Zoc18933l/qjKZeIcUTf5BcbWoH0WaU1+iCbrPZCQaWZDLNWuY9f
yTWbG+HD8/YrINp0gBxvntqiy5zZfjTkNs7r8xWfJF+LXxMoKsz+voBrg62l3jyzKvMPq37v3tPo
ut7BzfNvDnsIAttke43VPfO7nAJc7qkS8jXYdjfnkxIRvasDIa4oh3TYgqX/s40lyuoo8kUPckqM
06Q5ulYsG/nS1qriCkOA/I84u3zQvJ1YJoK41nqzfg88G4AFr+r0umL5a+gbkeD4W7Z0VYJcfzs9
zEWu0hTdPEyzs9/VdDvKTEBdSSUSjZSmtHvML6iN5YYhkUGhLXe0K5ZVmDnHXVtylCNQnRRE9x/8
k0e9YusmsKT5dExkwewEd0PJOpPWhHC/1ONTVeQ1NxYLOM/xkm4mexnmSdtvKANYrm8P4G7NhsOF
x3qswuIPTZU5haWnTqr1E3aQqydDHU3Qih1xSdspYOXDoISYk3ROM7Kgu57xRHmzFhZLmpEoe3Pu
4V0fPn+d3c6f71wT51Rg+PrUQYcBrs461vE85mphXplFs7Kwe75Nkd7t52htmAM9sIN8EKbpvVI/
q974xDRDxwNZ+L8PoHY/bzT+yWTeMoparclk3TuWtUrGVZuWWqAoNH8XXV/oBAncYeTBpyNH+aBK
cUhndwGWEMXG+EbS2W40UcVYddSWpBukQn1CCIwS3HVI16RSrNerYCMPHqz/iTiS5a0Wv+NkKOdT
9fIIONRYLqpk+AGpNX/07zPMW4KJj5PdGt1w5WEv2fGZFTPCKT9X0eeHM9L0OpfTX/BQ8catK2/n
30vCPNFVt769HU+C80USGW1E0HhTCy4YHMH4XhiPjeXxOPic/qI7uprl77BHXXh7uGL0Jwrzf2BE
3OEfdiei+7cPioyM29B7w932FfYXP5TqsUOLKN2cxFZSI4vGtpHj8+tut/DWXv0oLc6uaup13eDN
5Wt6CgCs2gJkJtbo+2+G801pYX9q025OGN+Tfl2KlSpV0Hf+505UXFKXcfiCBn5Z+6j6RE0PtcNY
/6OD1ngiL71aTAJR+KLlThSticPzqypmW0+eGUxJfmad4Ps6SSc2MwdO5vKE0hQUwyeg01rcnDSm
Cmv0BGjhXUkzxS3o1BsKf+5q1iUnlGq0aaVPO4pGDTK42MR2kX28xXWg/UEXUQ4C5rzd3V1fQain
//S1fTC9kPru8tv3oANNTR6tiqY/ch73oXSO79YxMMw7knk9oh4uN2SDFHCULVYNb+YEKTuzznTX
U9AhrtnEe705ftoXDWW2Z/5BDn2aC2BGVl5ECIZjWrCnEJvaH+lrPxXnKKPMVFwmY4s0/xjRKQdm
AodjXy9/HVdIFHDnU4wClq+0hwNvbn8LvzIKqBMvoDuIv1EG3JT+MnELgAVlK2YDKnkhLHHLDjP6
a3rSVt8bB5T1dV5FPDP35GCzwlovXu0ctfjdH867B8B7osz3LCoJK9T0PlCbV4KmNZ2v6fKo+6f1
yV/uB9Mp2mG9d8ZwfFkaICAm4/sdp7KqkoWnNR0sBN25CPxKvXQxp0idxIYh2Jqy/AP24p+c9SV2
8IHeLKddV5RHAvOSJ/7EUseVJevCzWw/PFtnshjN5V1MaVaO6FQbIlh/mDagLNOfCbVfu9GEs++Q
c5g7MBE7vg7KvENX5aQUgzeBbnhIoGk4aMXpWWRlE7tj892USPjkqmhf4Bhr3cdfFvJUtfcVZL4+
xwuZ2K7UG+dpAgMOnxISpecYQL51dcnvZjFEgLVedI7Tqwjn6i2q/M7kci6objlk5RvKEam/13FK
yc5My6rjxw/m7mmiLQ621YypA9Av5JH/lbo6UbNtQ7JppGEDjDPAt++lRYu7RSlfQCwo+TGxcPmN
Ub06GFZjDH2SUSWLaVx58fL3MTqoPdcf/2wU6UVVJ8tuvsxvTmJ8ANKL/TYupDsnGafiRYN1eVEc
1kMzEjfGSYWs2T1+G7xAgaEqWAB3XvifMWTrsK0HtmvNjAdPjTB0AcdekP+GGkyp1wOtnEp7I+Q3
k40M2CK9qrLUJb4JoYy1PAsPLKfB9Q+Laz0loPBAHVTKNswPJFKi9B/stHbtNEPT5oWCVT2Q3/KD
UmHWeESIYQnpNvmZUlDqiUcYMpCfa5C7WnPvmGPAdOTFXBg4tAXTvMn39n16OKVmgxy5QVdewaU+
NWbgcHKLCrZZHBVZHHv+zKU+9kumW8y7QJgEMCIUe0N87B/Axm0nVIb30hGa+NMvsyq659BAxeZU
AH714xOj4Zr3K3KJpkHgczJewxZHf/K5muzsR4h6W/3Uc9gyXiLxd5d/1q/Kdi7fuZ+KxMP6kBQv
vqVN5HcWAHdQBhGwrSgPpsqQDKkRPpedPDiNbViJknDKJ3DeXYpJECAMMi/fIyk5yUT+MI24uKw7
CZRahftsiM2NkaSCoDZhR5exrkvfS62b5UM7UZ89BSTxG+wgUgac6lcixfSoj0rJjE7dloPxKHo0
r6tQt+T42d8FE0imOpyhO9mb65KRD/VF8OEnY/7RFLr+qVRhATmDd+7rv65iGA9yvbzjFsGWTCYS
EbK110sYoHGUBuBcETZgTab9TiHckxXfPwghpVGf0VCK/AvVYQ1tRIwD63TWHO9auHKB7J9VrPo7
FRO5BSWs0MRKLpdvytxdv3+cv7ctJIBNG3UrsGdO/Kyn8P/NZEOopfmc7yMdxYLkAhWJPAKnOt+1
jOt0R88sHmLQqNkcKfexE/8cbsssIEKG1/PmbjHx3IAYgZBhW3wOmikwGqZdpt4F1+O7T+fGtp5c
Bh1cVc9t6tifyB5We5pIYyoSQRN3a4Jbe4Bdm8wASBDpERsEmEFqID9OlQraxklUQk1tV/idFn1M
roJm9NcsZISvYMRfQa4GQLRe5tz/ITxJOhOeigBIhFTq+3B+j+Lpob/koE0RPauVtzUud82xeXZu
Hq2c9TG5TlQbAY72KNRRb4wSwYLgPE5X03TWZ3oui+xYysQgPJWYfhaq/jEDp1YkRrJFSvGF/gUK
edZOs2gLgFuXV0NwtfY+UVxXxzuWlhlKaU7lTiq1Uw7wQX5EewqYHFiYtffKVIDEdL7edbz4++k/
nCKMYyr1euV7rHGyKqU6hJPW7uioCeOjrrHF4/yJT0i+JacZLLynHL2pxkF3eKMoNKmNi1Bh6Kam
I32JE2+/50LIewsvrBDGJq9S0I3ty7EmeYyqUi4O7fF/JbsJ3RJr7Kd2PzGJWinX+FLzWzr81e8G
cmGuLe85cNbe0vIL9HGxysj2a92JzUpmmL0pAaqtVcG1s+2OtVFmMpqkslT9MwSmpg76SpRKtfoU
/d2SztCy8u0yMAiha68J3nQvMScxnJY1CxZvi6naQUws7q6+6fFnBY/mfYvEW7eIpFrxU+CsTkIL
10GmtDIPF7GqnvdsL5qISVLVsefYa9S4eGvFsBgbkArXrqXYBb2ywtBSHo2gDEaa/X5meXDOZ3fH
XhioXkMKMF/9pU85eRNnydvXj2IAbf2ZC7gZXsL+kzho1GkzdoQdvsn6mb0hsr/pPncLSG/AfHGq
gDUzuiVxd+DFdpOuBwj5x3Mc8mxoVFCM2NOBrlMKdI/wyLg6Z0z5gQHNYmeqwM/fYUwCBTbwNtcJ
yFqfc+vpk6QS1Fl3F3z4k7bsky7Dycy78VZ+6n7bBl1EvAl5owZc8mtFOT9TNXoIUy8u+dyb+7fb
odtXqJRHwblmD4e6unBy42trf0ZsOFGxRYHIZkXY+QS3x0ZaGIqzwWtg3Dhdqv2HijdZ/jmt+85i
rW21fwoGsk4nUJd+YBlvtKcLc066OqeR4jz0DpnRODEJezKAkw6kmKUG3A3529/KIWa9RoK2VRfk
MsSfEsPTL8w2GOZQG+uenbABnBa6rWFolQusqpVsYvm90VfV727REN8CQECYSCWJygu8RImA6Wnb
V9zhfCcfY8AMS7ntrgVX9U9RA08MsWAkE61c7C8v7LSHIO7fbYwiCw79arSaQcBaX9LiBr8byzmU
Q37QIPs44yAoWSWPDkOWbYHFMYCX2rRDW6zkx4DDlrLAv5TQFmPEUDAOsEp1dmFRAjl9NKKChgBj
Oj2QPRCGHANtiRTEzdv2fENa1YPVrFCNUzZvYXiR1dG7LV5iXcLnICHDQYnOFPFF6CGfrhp/BmHq
mQi4QCBwjJZUZK2Ks5ZvzbVcN8avj2myVEOVZTYS1lfHUI/X1FMXuOHGYiaTFPzAsxzDELQXLPal
k9hqzhBedwAoUG2YplnBgNbkdRxfi+oB6mAbWF896bn1PXRP0SvShZACGlEyNCw9u5cjHUBs4cXU
NkBbeO6hJz3xW46AEfgsuIJXY5AMcNHlD0Iyzw2B8y2gio3qnjzrsxWTS0f1zLY4gd3LrpMZT5y2
SQRqFe1zYbxpYg3QCE0/ZMxN6l1C79IqC2kK8+IDUKpd29Ki8EO8J+yoYAhT8ru88J5pjIgDTN6v
W8IqXFL0Ea51W4FP1ex0ILy1A1ctgcXuC3A6+ebe1l6ERk0nJ5VjoUzEvC/Jc/NT7vrZwPmRANWe
b8SbJRPcNM31JFZPmEtKKREduBKC1logI8xTwKyUkJoyZ+oiqL/7CyXAO9FO07w3DRk2iPE/8Iec
lGd31X2JaedbiPrgqO7CJuhcZtG0698szmnFyw4zAA2OywOVVAfY0eCZNcMGAcl+MaBsLu97kYPf
etZ2VTrMiu6zDoyc1mA1vVtG7O84rHnOELgQKF/0EDiAhy6OxsHR2f3WfCPEk1dxsW23loAEiIzf
/HMvblvdqluoarG0ciU3NKOrH7YI8Q82ep0y5chsFMJFeRjVoMcDMQ+nkD19TFU/HnYi5/EkhffU
XqZ6IA8k3KPRpcThJCjmpOU7YyHMQbwNcCKf6aMCcdmOc3V1QsOv/dkY3Gp/+Vlh4jAYi2/FGgUj
sFYfZUC8rj1QKnUP2BDkMMSBLW1DizP41iSTItUXmMbVrHxSFIJLxznW5N0JNmnNpuG3G2mntB96
8AE9NYyobDYlLo53r72XgIiYkI1XFR3P67Z8pFYEIRwVKzvKNO/RF5PgZkq0GP/W6g8lVP6CcIoW
oAZ6ms1ICq/81XIKG1W5ipEkePnBlpu+ba1w18BosoYCU34/MBzelModnnNnt1jV7NcT4ASdiFmw
jwH6GwuwLJokmdAI6uj/uAB4Ihj+jGy1xRe5Nd3hGe4wYpa+VfbVZYC7hIrPUBZzkyD2lKLywRnX
BrKb89oMshfm39nRybQ6TEGk5mA3A8tZ9/9QuiEJdQuGBhRvsPNq3Pm49fWXIWp/sAa1llhrJqw2
DG2y6YNdcizrS3HGsY5acg9yz1CA043TKM/7D8t4m2LPQvmAPwZ0RNu5VM4V7J4SUP3DNidsdLwP
ZmgGIxZaUCndfkzRTE31Xd4/ahyh2JvFxo1zyM3BSPB56F6klGivJw2uNK/bucPmHdQzp3oRrrwR
LFS/OL0Ogt9AYC/6orAVCBcPDjbrOw/bAlmh9+rRzmstQE7fe7sEp0wObmoIwYs7RB5gxeZ2NVtv
8P80oGkqIUFtCUz4MNPM6LGR6ADDhKJqdSMFxCkS3vByIRCvxJ2alqVsotYHpRPf3ln1PEmes8Y8
V36n17EjqOUEv73nTcZR223wDNKhUm4pzhSPiIyKc6z9YwMI00oWjTu/+qC/MvFfL5xAbAuNcY21
qaLHHu9CZPp48KNY3zKse9yI/0ZHYb7Pd2y2lPtanhDVAfPszIGvGPsQnWJuGHM0l3L+zXCnSopn
IWe7PQa02AXOrOdeqyHjwLApfL2TEi6Nj1rkqf8NmmdiKOzoDujx0lYs2pMld0dRjE82fUdzdj1O
5aBtD+rJ2Asy+KMDV7QUiiBY00m6QCe5okmL6H24HWr3ft+zZmwOynKGqejl9mw4pV98xgcIHwar
kJ+d/G3u9/8U0hGp9sgi0w7Y5Wp4UcJROM/2UEA8M5iQ12ERARA1PPJUavLjJBWNu02Bn9UkzAV5
sJrUQ60PESzYn7T+ea1gGHcir4Q+xxVNaTr3sgega65gbtyi/Fi/UmaQnEhvy7WyPg4WZdzWJHyK
3mZ58CoESmnzuKbao5FKF3zl9EiNO9DWTtVAOBjGF7kEy7bOdJEBY6B4NOoupp81nEQ99OndRQrS
MXYm+uaH/JhIcBQhid8HPI9mbVbOAp0cbAsxr8rSx818cjLYfTIvhyJgcTHnTUOoOVZu1OC7su6j
W9Yhca2irX2LFgZAsRcB5pvLKw0PCj6LdgQNpXIBpsIBfo6jekQH3hELhd1TAFc9RzVVSpPRuGCZ
YBXjMbE6Sm2W123rlGUvyn7/4VL9fBIoHdTTsXwhTK1SER7hPCU7RDGza1qEJML4E5z9fzyoSrnc
ApUKLKGJfKkgrTx42EODGxU+CFWJAagGK+/XJSi+0rFkDo6xSVZFqq32kSOhIcBCJxQNXIvhl5vP
+tzcv1IEfTeFcpGuxx7SKnAWLN2PTOqGTq+x23nA5JViNT+LcxVwrKJShuO+/hJ1ZjoJXcj1gPpb
FNVykepuy+GLIIO864ckNB0Vjmt3OkI4mkLyrnE0IktrJ2mawxKyc0NkzkIkqkRrD5L8U11B611x
7UTWM5NN70XY8ijqr/Jvk01Khgvom8nukos2UwJTcvZ/7B4Y795pTlrZw8XBDhJV5ACDqrZDB3nQ
hS83E8I0vOjHkN0JZs9Yu8MzGhAgjdmCSzQy7e4GnArdhWsCggcEpmOaZ7Z3joj5jQcAoUMUB3EL
bqkMTxIKc6/vV0f7kAa/nki3yuBocVzcSX5Dop1gGInbApUKv7mVwutVV0LErfWI7xxnPOny+NBD
kfpQjifvhjFRby3rVncPIMvUpjoi6nzDRkvU+AOP3IJNivjPfpgZWAxhNkVDBbM9QhfA4bFDWTgf
xsITlDJ68k1FcvJ559YaWJTM1KF02bI3dA6adUT87nCtP+jRASajopCLp/pj6P28gwG2rMqunOUT
oJjPNxj8+s7XwIMg6msLZSMKp+bE6uy892x1TDZcTZY6gIgKl9YBJkqgeZxshmU9yM3xBaUQaaiO
/57J5QWyq6FXsOZSIUGEIMxK27PfXRs9IzokxCMIsq1InJ1qI2/uRvrNpGmBj/q5avzNkMrXJxFD
Pb3YUiPw7/j0K3MSWRS5KUwnXl/6gFkoq0JDyvY8fWA9/l9Vk7IIimcVByLeo/Ri/7EbHTqG7yL0
MEA9LGf3yOsgt4TxK1gV2Q0ROGqIlD1aZOYb2t7euijCva2vFnB7cmqpbr3FD/tEFJB1oM3TP7k8
CYzZF+8N3wW4jPL0GwVlyPo+fRewzHJjg7hMM3YagqIRDZloiwI7tATZayHaggdXRZr1l4enQnAl
V9ecVdn3R80t0RCv9m/PmSRHG80F+/HkD4wGKxWUeqo7RPzUeNe8S2YG61yQ3oW3T8EQUrt3eoq8
Yk7MGcCL6UX1nuP3WnvyciHkzhrBoN05OgOxUMC+q++wpNpw03O0lx7h3kqUMUivDCZ2wIdvAnra
x77xyk4FMN8XkFmLsr7Ah6571FqCfUaQ1m4gSPjE1qn0wok/rsyvEQ0/pG3BJCHS9Xz/2tz+TdP1
DA5oSCtKUSZiAJK8BDkQ8/f7rJvSWDmhSnLeh541r206jYR0/OMv1S3GYAAYIqumyePNjFMJnTRG
agYU2vXUN1LXXxhRuBpVE6M5h1r9BFjUijPGoLqj51DRV2d9yK2GQPyufy/vwZnnirKnpMhVMGBF
+EyU41Qt9s1b5jESfuuvGjtQfcvrzmZJvotwY75pcymTCE29koJjn8dMS/ljqTAsUZlQY13bwytK
5MXdDMiyc/bHJK7D/SrlRrubGY+VQStfmThRtWTMbE2MrKyoHJ2AQhM3+Nh5NURFNjWbw4630SwI
OONmpt34zxLLm7+g6nOAd6Tdu/AchECgbS7UPfMsbS6/GNa7GlucvL46TEoZIyKZdk0RS4ChW3Q1
SBmkbFTu79I2WY6kNB3CZ2NcOQdBf74t2c1KvZJITzeA29Qa6kSqhwanDJLx/b0tU1OudJjj3E1h
kq7QevEdQqfvP6GluYIm8VWA8+UGQ6Tafc0oVYce3hCYyl4e+sBldmVuCTwgofcOcIooMdMcKfNi
w8asEuyVkSnPWWCw9b+OmAqwrQft30mYv+TpBBx7QWz9LJ4cxkDv58TDw/nAIAcrWciWDE66J87u
Hsevr041MXyxA9+vpiWuLE1mibWC1GEFXa20hQkBRZ9x2reTU5XVuhkAAabkAR9HbqUMQm9dPyfq
oAS3lCz0PlLslLKJalID+oWCT+ldHL10m1d+Qk46awnPeBQYFwrAp8cpyDK+h4qXmjvwgYEpKSz0
Pf3Lqq2XdPcgiWpUC+tObkozBEGa/oNoBDQRrqUBEHJF3DYUnXxMw1J8pP1PSdlHfsWI/yISeAny
7pHcKSfkLhE2BZbxv4Sxsw5+GsjR+kwG4doxmvGF+PdsdprxliKRbjdzDsfawhpxidmRoGxyjL7J
O40N9Cd0NeufE1S6K8uJDFCN1f5Os8vJM1uDWGGo9uU781E3ffTjk4KH2aZqgTOLPIEqtygoa3SB
/GmCCNcZr2ylDwGUUW7OIqzNs5OklgIiVtW4KJ4VcJlOD7ZnrYAuQYc4lZqiXxZ/6UTymKZ60MQS
ohjwzWPElP0rz1iqr85lmIosL6ToLNCMW8UMLR089CtLFQuEqLpfiKV7eHOBFWSyWR8rg3Az1cwg
ysKNJoRPukh0V+FW5dP7xhXY8wP9O/2N8356k8i9nqaXEfBEbmbdIpRl0jKBj4FVAUWbocrDboGI
mz3coa5bBqPr/MgBtM77PhecHpTkYjyFyAs8oDEsm+Y/pEY041xHqxoNSGZugtgFs1uyagf738u2
3UZnDPwALfZJ9X8VU4nBB58NspCZ4YIbdoPrjKR4UL7WltiwuxnNRHyTOFA7S1pHCSPIbiVNj6dv
SgSo8NiO2fVKR5QX83g1ChLSiic7v9NpzXe7ODh1M0mWkuzr/sAL/EbtwGalHh8X7/1IaHRKqLgy
LThIAbyBCUROms7STNRgbuOQbcyLcjc3UpggiCC4QL98Tt2YnaDWyWgskQAKSPrZi5TBZGQoZKBV
xXO7OAJciYBdmCj3qnd+LjLzLIEFTdETQbtA4HCpORtpfG8c6ciqj1FP/wCyqNbMTBra1R3IfAjw
+m7hPbCFxgyBWmf30GdYhx03I+QPLX/XkZ6KgcaTtBQ3+PT6iX/qvRUKxCLxo4eYGVKnYL7j5M09
6aYuX5IzztmjLexLvXvMfNf+M6cltKj/uova2o51umsTEYzLhiDReoYOc6o/WONPKmrFx9apCeF8
IYDY2bh7XfGoAumSVl3HWBXpkXqMMWBx6ujHm26VmViRf5gUX+6cAHEXXp087hk5G3qhToWVQdTr
sky8PwT0vJM3PfZkFQZjQVRrbNUPO/jjsTckPnW4SymcYn2Yq539RGk1rt+Y2HlUFDksHgvzC4CB
5ieMCkEh2UCcd+aLyGoZIIg4GQllDLgacb2fl2u9IGfaMsIYvKY2scxMDwFEPXXOia1CmEB5ZcF3
3fkGiGiNRI+GQxeJCtTz1FWrkzrEh9qluddNQ9Hf5LmyC9shPNRmuWOt3kI0MRoS+s5mqFMJJRz0
lOSQ6CcXVoOCC19KLSdqESOZ8qgk7FDQ47euBUo2gNBy4HTViD9hjpI0mi/RxxS0HWpE+A5JFPzQ
+rtTGmy1yburYSdyMNnEiU74mmj8klePX+5GhjrpMtyePGAJp03RbBjcUDEgNvQly18Io2TiHWgw
K0Kvdss10XxT7PKJNuEMaYFZAZ42dFaciH96pJ2jwAOcvLpTPnc5V0dM/iTOHnb8o0FQFnPzTPZr
wb5pk76hg6duYbegX+AuP8/np6Vf8hNjI9f7upNg66bx59msjcfi9DJv55yy4qSCp9d3tRLCb7nu
aohNjNezA9C/BIwvRVX8J7slJOGWbRqgx9IYzqvS8hshbnNkjhlsx5XSkGWV3LZhhl9xyyJNDAeQ
Tt7E9Kr4Ld+aszEpRSe1U7dEVNw6UZhnraGc3aqax8K2hRDsCg0QZzjdEeJzGKLLQERY3pl2B7Dl
mDdHfQistV4tBnGM9NAUp5ZCzxN3d3JRDuzjGc1Wjy5PS0zsqF8KF9h5V9Eata6ny57liH9mKViB
meJ685/dTkALMQe+vx0nFJn19Hd9DejzWR8blmhVOpBcEgwT8iDXfTlTpHnqAjMrZnXvRt/e07rM
Lgz2PGMaJdggyjLvrnTj9miAd8I524qefeaSxmvhajBXLRxg8Z047FfXtdOaOdFCPVDqq/R2OqoC
1BgXoJiwx/nsYPHBFH1M6F6SmLJaIs3/XATkin63rHt80DzsglPEI2TFoCAq2HBQXTDf9ETT5j8o
2L97cWToYYjFyu6fz+A7Att2QUOeF84Cak6MdwMEizRD31RAQb2FEHkETf2unYgY+sPt7zl3CS9O
Cw8XRV7ZH+7BJJt4SFUFFithuqEk6412Jc68GN6EWdbWu02AzkpZM4E2cdFuhAbNyGBOat7+AVZI
KKRwCKZ/B2kGODuC2gSyCUrgAv/itjCn9lPKSp7dFCfQz54X+2/GZIgZER0ll1znj7Ps8yx2mStm
GYvShf2CVF+Un/zJvrz0s7xZc5N3r50ZKhoQ3P9b4CH4mdnnIAP+j5IMRTtsV9wniEhZj0WH6UYD
ATcACurnCyGJOynkLRA2x0LgpE4TCKu+ss5Q9PdPBN07Irbb/Xt5UQgErNmJnlt+DDRaiqDaGaTV
2e6aPJRE5JSPP/J/O77y74C1cFRxbl6yzkdLIWRQGbX3cyulZJ3YaxFGu/qeBuLcLVjsNeyDBwfj
WK0vBRqBYxT13iIPTGCuzqNtOTA/D47Ay/ZQOHW08UjoQvFPi2312v1OCJwanAmqqhLLVe0yUHtW
IztfQn2v/37f2f7gwJn4j9MV4Jx7AvY5UQQiBfInNrDw6MHn7A3mcgAGD30fStHPJyHhbCfWBTJX
zLLdLFNVB+upu2vZp8/PxhpC/5HBNaA73MjgPynRdqlu5W6zIhcqI/4OEjYryF/etraaReCG3gPI
XcLSYqeMn2qsVRgFTL2taudjqzPEHj50KAwngs4H7G1jfB8y3PEpnUWxzrfgZz9UvJnfTafKqJco
tNVVxwmXyu9yemIaoWfhDbru21mrTO9y/gxnrvAXrfYbYrALIcz1uro/4mZZHhl2+Mgerq6y1USH
twYTPp7ZW4QE1KAbtCtDpBkUPY0vMr6+32iMa2PEEss0mK2M+Teg5RvWuJcYI6ioWp1jE84yr14u
m/QZWKoGFfPgt+l4CMqsE0m/uYzX1J49Z3t25ptkxLyTR1ZsYzXcmsxZ015fIJ5cHPGcFbGiJRqB
ProqA656XRzkBWMU1g4i8xRLO9kfNY0KnnDGX8a+PPFAyy7+L29I6o/8yeHaP/x5jDaSrulJ2RDK
2yYNvwpAKD74sRTw3rxLLJuv9Mn35QRxFacCdtGefDmhQ577QFBxELn3ONF+Sfn3oaE4veQpHGrH
MbZqRPEquHEQztGbcjC0Et77/dWMFo6E3oVEauSBEQC6Iw1g9ju+DY4n4rjBwFNK/sOBGNotj2iV
+QGP+i535WoqPRI/iW5hOWLWkb6ZoYOjmTtYi5X4+RQEB/7j4ZuoJ/RwfksbSAI9/FuIPBLeBBc4
Gcvg7mXtHwGyA+2uSTzfSwUV46uvKYKnFKlcpPTQUD5XF9h6YoRQP4IJwTnnSX9mYYnvOaQpRB48
qfYEPmq0MWkyYMRaBxJaTQgaeqHHdvoUnD/lahtGRn2aefKskXyymToxnT5CU33QYB6lY2J39yrn
FbiYBcRwHfErsokvAeeu8o/rtMrXDJ4eubgadKZKtYx2gK418umuFgEJU7ceHDLv3VX9ggwukY31
Oe0m+nvOKdVKf+mEGuMFjoWFruwbhCbHMzcTO05dQN+ooPyCjCbEhgsAGiA0f5KaAvIHLu0BvSCL
WlNmPmA8Z4k7t4Do9LiIw32ryFePAwobA6XgXpJbjLRb0gsWG/M01v8pqSyjXCd6wkYxP3Yuujg3
+smUqMqQRbhp9zy5pX1VFvRu/9dCO+IPMJ5AtoBcBKLftzAd8Fc2x9GzUiut/lzlCIeXK94zZUpR
uYh9ZCPGo2xQ68WauaKxvcgc089vGHvgL1wSGtsXDQaHSKF0J5Ow55F7LrOjhs9Djb3uz2zUNzJ1
C0tgYwSJ3nA0tRiiSQe1pt3QF373iCAAzRZMcIRIwHqFeJ68XNw7UDuATV4GrMvideP7KlD7qwCg
dpmfsPxkTXTmbu7ZOqoeT9oPmCfjBkX1mFWaLV4YP7ANJyQE+f+I4Httou30Gigu7wLMAuSETkn3
QT2jusMWIBHal2Jt2OoeWI41baIBJFbQmCjEgNFESwqjtNtcAfBsrd5x8tMgwC1TeUQuTixWFXTe
MaIELEWbcDq3QTcKPy6wou882Cg6yGsZUTqRkcLOhlH5SMsZ2t6zcyEISiNPsG6sY0cFAO+x1go3
ueAIZDPl8tCjVPfcvbBq3aK3QfSB12HSFyXYyJWOUjD1mlBpSHMft7jg/XoDlDxzhqASXxYtFftH
6fBKI9zhBFJ707bp8+l6ODyOA3+JMeutr3TeDmJBJ3YZD3QyL5rbKy/Jpqs0/7We+N09zPH4BLxq
UTiMmTt7cp2z40EMvHD9bQ7eY4yk3IeD3Ad8aFbpFeWVCD9axQCZGTEcflYc8C7o1irL292ojRym
u13sJWsCYHlayYDliGQyoUzWQ2IVpFU9MKUU5yE56pIgCHoXe4Yo7J5jFzwaWTiimTYLbWie6ZIa
aWnBnpSrL+N+LzhrV3A6avjPx5hDDsHpcZlS/SDvvAdfKsJ84oiibpIHp+2xzgUfsTsNLOKYAKs5
HayQDKFZzz66uASbT/eFR8pHptAU1GopUu3bPyKpWZ6hG76OpEYoA3j5sqtT90P6GtxMdK7Xqqde
41EKQTtWLeuLRMnTuvbNX6zjoRd8vzP8G9Uh/+vKEBqNkv+S5UA6+a9hWS/1T0zyH3/OVWcdU7uU
cfgWLOEUhrtvam3qieePXqOLr7H3TstNwJWZH85oTy/VhIXI4V/Ysh7ATkgJKU4GsMrsXTDzsyXQ
TTzkHv+ocxmMBWfealI/yVkW/e8Zg+bbXJXp/tfQTQZmHzjPSGpb4oYs1/72sfuRB1+buf3HK5tR
No5chxTd+kDUaNegpj8rzsgzg1kTTM3RNgufadjTSsoaM01qGeBYJtXjt0wXFSwgeVFntso/sDLg
GP2gS7Fnbbb4iU0JOx4YxXhKFn2JFtAUz7Tg0MwMahzHDxsQknINef+Ea5H7rQ6l/6QaPR9FxIXW
yTIZWcIAEnr0M4pEZO54nIErNEzWB/Qm1/fqHtZU8Wh4bPm0Plb57VlcUGQb6PdOi+/n4VEU64/Q
WdzzWK6AS6XZxnRdHnN31E9jN8kCz+0JaRzl2rfl9qoXTW4RqY9LiyT64q4PEXb9bdcOny7TQDl1
4mODqHZ0XUyazEkcrpoN4SU8WVilrxHIrhCdf0lxVWCBnhl7HsCeQRjk6CuOmEKM1UjZSh1b+rpA
jCQjKeOOPxb9MdttUjstUznHZsi1tcavHxBom1P3+3YNncBv8vbaRFvCdJLeuQp6LtynQnkFLBL5
b/p9hSMFwrDBSNRXt17l3F+S88PrMuTU/eDKcl4Qh20SvIHk+1ZMMuw4pIulzO6etZSOcIVcpOva
zL7wOKZBn2Ljk7zpDGOeoRYkreukIuQQzV3H90tZ866vgq22X6jY5o8pzd08O9EkWTSgYD5f+rrj
eBDXYb5MTWB/dcZym3i1bMVUJxW4otQMAQNLeDfvSUr2+nCRevIqEw8BYxiGMmykH2qWkVur9Olh
LhGNJbZvnJM3eROlp+LXt8w3eVVlUP6LAyXTAtYJWN/svunACYN2uNHYMsZ1PEHiRPYo0HjRzJG7
Q614kAcNdErPJjgat3GMElKqOMh9irsD0mN3pimSqay8Kv3T1zE5ehl6CuDiQ5C31ux5cLayVKKr
fVMUZc3uBatX3/m316ng2+J8SuAsCqbHv6Cdsf0nVioaXeOh27a5IGXy6QN0u3UkZ2r3cPI4TI/O
igX+eTNPkHX6C9s38lPfjFTeqVTumEzpEfzrLSltncdyNBgQd6ZbJ8/JabU6+9vY0FKR/cq2YRLJ
5hKiMrmYMRo7nl5evH6QByabCFS7G4qC1EL+aLmkNMux8Tl1zPhZhUfxDgVeTAudFhd34U7/V0Xu
gynt9lkHFYd0Pg5OmaCpuv6SCHpEjtSc1REvFlzpxWj9Yi3fmA2R8kwel8w5MpZfU5Y1O+0WdlWB
lPUEfPQg2+ZYtTqW7S0/5Hx74dOVrPz6i7AFGESFnUBWKqc/sl5FGhWNN9cBgnBEy/VFiH8SnCm/
5B+U0B97wGG2AoACj3mMlp52crMh2dTUNU8M1eQMD7uYdcUx5V3o/Rqr9ys2ZxwVUnBDNPJID9px
PrfetdboPpdHZgWdP04MsGJDTHRh2hBzxtf8RG34rOHysoCESUIP0sK3v0Z4Hg5A6W0QUP7rbOJo
9AwONDlBKG4VNviSJv3QwXsm/T9g+cHGsXA9jiwOhr7nWwNAM0g8g1jA2pz+b5i4gvSZpWwO3xbz
2hCY4aWQgBTPISmfYsNggJBINjrznk6mwFIytSr2A1gtkpGouMy/y9JBVblLoov6YmU905TQokZX
3lz9uuYwUHF6FMt87z4icQ5fPMiE9HOIICZWYniwxgLakRpaU/gKavA3SzL7E4YVlnmLumBpFheU
DaG3fglHDEc4u/irvqvNBxVHmU7f/+bodWYLKU2AJbQoiU2cGlEbrGz226fqiII2dtRsImo0wWnx
Y7WWoxwOak79Y4w/Gx3oez3yM/Tc2VwbWD1hG90DuXxf3My5+oGzDMOp0mh8zSqqKk4JKHOA8H4m
c2lAE2YtcFxoonWIbwjJZBcIUDsKfRq8loCMUFMTAcJnSJfGXUDSK5C/8EjBVDXJ1E4yXZ+TLqiU
PGflNRF2LYDFAZ30MuPO9VjmUl+p/EQy0tVlflRXHBjr2L063+0rdIdGl7urLpcVKy6nskyuH+pi
5edkBm/Zl4zDcxhnWuK14bkUHQ3EyYTsnA55q/UTflwvXUM7/gJlvPy9gKCozPdWykGqhZyaNWT7
xRS+Za9TKbEOXLVB1fPPa5+sqnpCXVhg9YUNqn/dLnp9MhbruBzEFLSvVe0eapeK486wzjNX49Y6
tgqekveWcCmCBogn15IDxj/qgQzzGhAWx2onQsNDRt0IHCE7hkSq8CZR9kDOub1Y2xVEbiJ30GXJ
0VKffHbtStydKqu53P0ifZ6Gg+K/Sxe1mqKi5njwu4T4bWC3bheycSrxlb6Lsuxft04JTyQ5pQbi
tHYm6pA4WQtqi+QPohYt5zpLIefP9eBsYzzZ7R/kpjDQKgJvYLf7H1oW7g01RRYuTqDp7I66Fjuz
RZyv2escnUQG7xoIarSGcHkDS81K+9MFEYhZHl3XPQlEE8sTSROvwuBMZoAqtsvI40zOf/YzCTaF
NNUIu+MB4Wcaa3SXXUQJh2IDvuqyTo4Y2NcCcJHgGW/BoBUJ9jerQvWD0v8t5MMs/chcD47Au53t
D2HGYZ+WVcffBfVLUrlam+tFGLti5bZRLfKHUHDe5MuUuym33ULXBJTdQppFwW1xG9QdivZlFwhr
2h9tQtGDA7XCtJenE4ZXmWY+l1OXY6qOqYR9v+XTor7LJDpMYkRwEW1CZyx3DwyaykzNTpvz4R4a
wAr7JsAfVT4APB4evxRD5wO/1YAOiRClv8KNfr2cOl4qSBMZ3mgLESDsmuEZY7k5rd05FQywfEId
1q4trjuwHdCgSryo4GjATAx+mMI8cfibN1NgDfCRjUQznEBrpCa8DCp9HpKbQFbZ2ZpWqY+t43vP
nOq7Cr84a+H7UF0jOTR6HmuyxZ562C2Fqat2swnXQ8HESz8lCLM8Z1yXbCIb8XpWh1Z8Z294iMbH
YPgUzvSLPZ4rGYxY3mK+NRhkUd2olSmiL9eUb+nxnTWRz1lbrEY4oW12ZtrOcuVAJz58g7+cO8OS
jkktPkjVpsSJDSOE8te6LJmTsSuJRUpGujXTpxxRziHoiczRn+4Cbk7x2Sn6Tx0+cm4EuMjITGAg
VqrULRNDJTdhpIxJVSv/LNp9bAFtvKI5xaH1wFB36g5Ui4aHYWwhqNl89um+ZQDyGowuFBApUs9w
TQOyZu0Dv2fOohZEq9au3uGoZvFUW9Qu262cAvA/pZAnY7kEAMkeGXkyptuMFn93T2OxYNw8DEmn
uAeR1LjTzpNFwlGIRYItDpxqCBk3MvnVONI9v4xXc8seZ7OyYt8XKWjrUco/OJNj/WjuPU6IvAeQ
0nyzDfITViG/Ygb0iX/HmalXIaFcWEfP97omiEcanPUKUE/DbhjDU1ZfGh78ENUlcD8l1RxNqd3s
jMOAtSNfNdu+bREzZDzOSbOhGDoqYn8w/BTamgTjcQflWE/hHgKyuZLg+TLEgZw7jrVRJV7anYy3
WVgK20ns8NScJfuK+Ffxxi8lZ03nswCkWdynuXFnWxsbzikHoRGWWK5/qmWHIH6x3Wc3hgWj6BRO
haaFMTYQUn4aPa5HlJU1igMWWbcT4Iut+xM75a1eb+i/WK/4KfTfXwWz9kPPgRFWW1FUMfk/dAsT
15RgryPOiIByRfCSxmrKK5pNlrwRYbe2Mhc4OwNi1rHZQPEO6s12LprzZ0YZlJ4U6ZRZ/qxnm+sn
i8QSuz6lNd8qAZOU+6yHxuGD74J3rkPh1LKgYgsnongZjZkdSu3zYPeYNccehD3CSf6K8UGqBjWF
Eh/y25cM/B0z1BnNn4v102ZtKMD3hacanC0drpnFlOmGbVri7RdwfYX+xa33Wf29jlJutP0prxx3
BGSNKjEd+LphyFRVIlxmG4xj+umOFhoeu0PnpMxJIV/GsFZ0d5Em+vargrHTSV/bJ9cash1LioJZ
kIR4hpNfDLXs6FATY8ZEg2YpMSJ4MWuGUNtYa5W/nXCKXqwYq9is+oq6aXUXPhwO/UkQq9U1qn3H
q4m8BChOVomXjoAvPS3twuuJHiflp0XbGLnJPKA46XM9CoGcAFUOLvINY51Ltq8PooXFfh3eKeYt
9J/zqCiD1mM6gc523ii9iPal8PT34/ezjdoaJ39HQwRN719XYXpr4AOJw5IPIbj5f1RWLDes7khL
ttFhWUQJvbYCsKK715v1gUgfN6KtWjpI35F3Gb/La/llSCZmzg4yXa5vzprnyqynp4JTp/51eQHk
maB8LFYsDZmgMSh7oN85Fc9Wk5b0FJB0pwv+qkVFbIFms5cxz896j4TurDlUcLcRxDLuZTLhEWl5
MXFst8FLmJTcOZKcJBwd90apYjaqWNU8LS/1pInpsSlMB45JFanFEysAc4P/i5fc/QsUZ2fXr0K1
TQaCCOrcz6QbvpIqW+ZX8mLnDt7OabZeh5InjyG3oCsRVWZvM8nnNDZlBfTvwGvsUAPLcPjJM2zg
hsa3cJe2H6BbasKD/gV+BtD4Engk8XW8zp+UW/A4yNAycWO10mQLnxMY6VVLwqWxjCI0wXLe9N0i
dhvB1CxcZRIaTzenPuOnN2YVDsME3IC5MHmzxgffZb6i4/hriqzYhZzkb3mahk3MNjhi/gfcryoX
N1d7kbmxkNQGAGR8JspnPYW9XC1yGKq9u5x/EP3jVUihwu5O7YxV/Iohfs9aWLhHEUZ7h2KzAHmY
b5XAKd7gRgACFZu+uZMD0ebGMXj2/F4HzbatlF6vUwS8+F/ondMTWDfO+lUcY0WxGDq7JUGIXNDh
AUDvhTUOBlKYNtpHEp5n+8llyoFtIMDtXMN3BpbcJoleSvZ1LVc/DdFiLNLIiymeY6JuLybBltiD
MrB9JZDqwGbEz2LDYeedvOWE81nFgOAwcWIdiJ50mUVv55EZYGshg/JqNZjL+74tmHOQWh1UOFx+
n3Kc+/MZ4TxTtqIUnIORf6/i2RDFzx3R/4uO8IZzBDX45yEYweraFQQZ9XGMPY6dlA10rccfsHl4
UzuKOKTcsqw+u+100gl2k7jCYfHE4B1LhfTw4fdgwAyXPleR0K7cLyVvDx15sHOrxifb8KPgj4zt
AnUrSlBQrrULqk/qsha5Gv1HcH1AF5KMVNvK7eYXJTXt4pv5/68Eirzr5JVTB/HGCNphiKlcRNX+
yYqD5RKdkrmOg6AyjM58b1ct3hPbRSo3SCtndSXY/yP5GZtXJ2E9S/lXIMyra+ubBFWxTA+M+0gg
Yk7wxYg3XyHbinB8uspqCgT7FWgUqkgTrKANciGK7h+J328wPg7iuCwBXZvlq3T3xYLlu/B8Hml/
JnVizqkwAhzxLkq/GTIVZ1Xnss+5igoYVu3s00Zl6t7gbBkqijwwD1+le+0RvzN3o8Aez+w7a5ce
KXa+9EZ2JD1VLTiExWqjFtssreE19XL32TLLC7ZK2P79srvNbH7bY3iW0Y2Gt09pUH2fg2RciIx3
c0lKb2MehI5+lpQ3ChUqgFxHzNbLpqSWZp0DyGckV3LGnpUpH/uI13a2XINMHf9XE3+VoEYJOsLb
59tY61EVg0T/4pzUO6jvFB9+Xf/AI3stKOeksQ/3CD5QMifMIwJeOkcGwXH4x0jp7OKvHDEwu9ou
zVWmNz1b9UmIyK5r3tg9w6uG9t/H5DNqFY8MF6s81vt9N+TFAuZqoU/cRAgVeJLLOhQAoPW2sCSb
knnVCL+doQ/ZtBNr5G16JgTrlQV3SfwOEsZ9jNqmlSK8TmtzH088lpba+4HoJcPq6URMb2LtTkE8
xhWnEz7UHscEed1rkH5me8UYJ197gTJ+l8FhEJV9M5N1BsHYCjkHroZeSEtrhpDb45v54wMYW959
pgaixnKERwbwg/aBKz6Uzlye/n1VzSeUwY1G2ooVSdRY1U4s4+iSETTpcrOE4zazVE+55OCGm/sk
QJGDbpqPBMIJHeI45ea3+ge96wQXnw6gTbzzMNZzt6dA0DDY6y9vi6TYANKQaGHnslvpEv9y/jXr
GonSbQAAR6YFVPZ5hxOdAh26IYjWvDTTWX2ssnNugtlC9B2A88B9oIevPsfugIZ3vR8mpSNIZvzP
SjO4mMDeX7FOc0gu90obzW/bB8vvClWLN2O7LoHE8vNJj5PTQj48EFQcKoWtIqafjQs76drzuMyG
J4l7VQLxAQ0CblE1DYdGiD9wm8RP6mvqDiAEL8ASP1KgrCg8hk34sV8oH5ey5AuOABF1XIt4kBqp
UD1eAzoHYMURETawAwWYJEJOUwH3mDmZlfXqw0PZdWADLDft274gp+JmBoHAonWf0y+vlzNe9zo1
524a6H86PTM/nNS45lO7fOnLNloyQt+dHAdm0Ozx7kcqmpadHiUt8b64Qo6DOVWlcHMGm4/TLgY0
u2Lr2yxy/nphXG52lMgsYFu4xwEI9zqhTbjLNxf9tekmjhX8EiaxIIr+s8dSAZjCmcN8KmJK/0NR
RNiajyKRtOjsFTdNTJ7cKW1gJeIuS+NtDxl5KVrbvSHiFhHOUAbMPuF5fiorKryfX+qrauQJ8+xd
JCTfXheeKWA1iIYNUYhDWPr9z1MvZM68eyuMR3BqXQfXQx1uhg9+QCnRtsb+ELcY1F0SqJAU0M92
OFMeX6rMOWRxdmbgoSqMRvkYKu1yDdseIdfBUmhwAZjwd543lsA3cvnS8AtS3ScIRmj+DyERvH3K
cAAacAMgPuH+x8tYOq/PZG8imz/qaVjOJfC3PM8jhCLpaRK8hC6rFA3KW4hpRZ/Rzlf+3e58FLxQ
eIGKuegg8Fh94yWZFUgV+KbM38AUv8TJBoVAwidhRaR5ioqgZ7OroLjIiwc7HWlV3LgrV2cnvjj7
Ogn/MXrU9VLFFDT5zl1+HngTSZG6SwMlEbXGmdjbfnpr6ySEu3RHETBBA22MpUkWLTfELohsJxcl
JSy86MGAqeOi6FJwzf3cJCpHS9l3Wy0JgeeRa97B2StFGPRyCjhOlnIAX0KTCxdyxCHsSzgf17/H
yLYIb/ZXLYzjtTcUN8nLUwQ5prDeL4mXX5BYYgy7rm49ou35jChvRy5y3UtYX/+hwMngVVOQsrmh
UzxoQw4/V3U8veg9641/wLA0/x7PHVUZDNtacaosT5FOCTxzQo3Wj4nghMHgmz6U9nD2bG59BzJb
VxVEXeP1+vYugKT2vJXhcSsb3lr1TkRU1ve85g+LRF1ruVsYQnQSV1+0Qgo2INT9OxRWVOdSnndq
iRa9csgd0knGaL/fVy1diLkMbeOmlgXXRUSWFAXUu1bFL2NwB7oQPTwO/q8tb7qFikZ+1SCv2E71
pc7Va6vRmkhcPtzwzTVDfL+qjxm6oOEjmskhR0ngd4GVNia4Nmpxqcp03LPfipYg/Y5qMHkQrshV
1pHssmAi9LyIlG6EL7Z2CUNRQid6RByeMoHOtlYo4tImnUlfNnZmTDtpDpWa9C9PIdOGg/Mm9Fg6
e2V1l3Zl5pnsEZZDFqmzTXrGnOPsqIl/9vglszSXiCexKDlBABlJDvlO60KRVZQFYderKn8KgPrU
vU0pRj2sP0XcONkgGJRpKZj/BJDwGwET1bJW3rSAH1TWbibWCjz9UCR349uUe2SM6Det/BFajame
TXqVYJXG5t+EeBpkgH/tA9wa6jMdqdD4TojiXsyX+ZjJTiYfFl71nhbz2kxcfsWrw2BkQ4NIxAAb
oCVPb3K6dp10pFQkr3Bu79tqZStJtuZRUOcbG47pyVcKEKn39FF1meH4hRArf3upQ/C9/1YmUCkH
fGmmGQ2353Rp2aIutD5CChgorYpQvRMKsn1nOLzFWG0VqsbHa4ugM1mc8fEXWw9uGf6DgyWZxJNT
qd8qfDjfFXwuqwsppPYX1UCxExznIHf1ui6XDif5Gea+k/MsjauY13cfko5n97BiMhcXjg5eL7Sz
NR3XYE3o130l28bSmvj31DERY5Hb8F3690VjjTdFFWnN3oTKZ/D2irv/F0b965cD5AxtG6HJNmYo
GTrpoej3+HAKhbqxhxAfL+CT9ekNVjW4nyRG8YJc+tdzMBaF4RgVPXuzBQUAYZiwV2vG54NFDACs
wx8qTDVL7pP0kgCKWYnf+RKWWlRfGfOTrA8Hvqo6j1k2fwT6++ZpZvzhzzIsp1EmACEnYX+w2tCx
gZqDvjwKyZTltkN8SoKQtHVhahpfDIaEM5b0/62PUfNkcXjfleYJu2bJn0BMnaZAMamVYGMg8zO6
wwXOD6VfddexpzFXMZ6NYp8hko/EYteFrUXqcu+AHP9S9jI13UJ5uMS+4uHcCboQd+4QY4pM6Tpr
tnT5mHXpuMTKc2pdrwDw9ct8nOVvgXMqSPe29G6aNK3E3h17x4Jv3zrUqqnRcoHfqnhakia4nPqi
xX2k7GjaOfFx+ajtxXg2+2M1bVlbt/DnFI+jMFklUMIXZ9hHXTojMbAWtxC4YLvQohGh2hI60qzC
DJjzQodPBCE0MZp4zcoKhtT11QxODkZJ0Tf9MwiQu1d8bocani36LLSKnTaUsUW/DmUr89OuWLgh
lz7Otur6XooHO02eLaHzf99a+yaXiY0JQfJO0FXtmnVeiUUckdogd/BWI4E1u3yQU6cDSNqJV+5J
iS0pga++XczSj6f1PMCQTvuvcojHcyKo7dVulHc9mGZeHY9kiacTI9e6eOvsy3DIZGm3VNENdOs1
Lbp+QSdBaFL9+1iutEwZ0+8EtQmfvzU1E2kqGLGlaUXOtJ5pnJagl/9Gl7h7YxiE7KcCCv/dUxS9
+LSI8l8/7THcTs9dGaTe8S9REJceTC6Grd3c5nt+fWkvvfJWDKz8upRe6rNeC+EYUTdrRkvgjKZ0
8kDBNVgqfdwDTrS/sXAFmdDA8zM5bboE48HngM/5ifxZtJhCLUq5WGNjwnxY0NIXU8gAgTAG20a1
n2Lfs9TNhs+BKdnrHN/NrTeDUJGUGNQVFeU3uyVi0JLQ/scm/BL96b3FhKclMNaPJmfmrWOSw6kT
PmpzhuZGzo4N6EEBP1EmFAuQl3jLAne7U50YiZRmcmY7gSCuiKDZEQIgKD7XBN/ZJ4GPbrb3g2mb
Tjm3CeouU2fVl+o/ZyqAQI6zgwhozF0xnXkHMQjy1JzkhMeSDMe37iVa6qnjB9GlTCN/nKR6TMap
GZ6HfHn10fHERniEWoxyLl67DJLOP/ZIO729xvb03DGtJiDbCUFCahMkgNoRTMMvoTQVk5sqSSUK
OQbLrCHqa/q4PLRE8iY0TZEij6/Exn9sKQVFq9FRUXhLRbq9Ss4MV4NmPD+fUj4vXYuK4o/Qbqgg
KRnU9R6T2Sgh2NeTIhPqLm5HdJBD1thxUTkSLKBzXnIx+MYtZU26Mt/JXExV8z0U/7rB/jUxVcB1
EWuIwOMphb1c15PFY+odeic5bdwItCH6rcE3tVQMeesY3/hPSeRe5LneCXJ6XqQuz5CFNxeejvZp
TFXCrVvysGZsVe1HsOu1WBGNbMbztgvu2vUOg4V5MQql+tiIrWANNy6rn9TuzwirQJWkGQZuVk0/
ouYd3bqhX2U86ow62TNwFZFUs9AXBAsVOJOmmDR+/O0yzd2vAJ+d/62KBCienyTpFuPDb4lDc/LA
wlpscFS7ITuVJVT9N5bctyyOB9of08J/++ndPGrMEjoB2EdtXLzv/pAbbNbud1p56rVonuCDeI8P
QlWj1Jbzc6QCUYVoai5nxqcSujjjuUlMuWYM/VUm6XhqwAsTr1y746f44ecMRYr/3l4wd0z7HXCN
UwLWtrxGSCqgr0ZxmgBlswVTG1W9yjQsIV7oM8xcr2OTExZ9ffoP+t7VPYBzOAX0sPylhnBAUold
xCY/8VgerLX95QXq5IEFW74Sd/EZ6Ot/xfZ2dVfGV/PI7WSbzEMKd3fYTq1xyMQrYYBURR5u4Yuw
Zzv5wytb+994rdpGTGMXvP07fckJFB0AaMEC6Dkvs+Ekx2l6KP95hyOBpq63lUKnwvLUyZFZIUXO
lF8KQRei8CkRoTZpscyLuSbr4Y3/XSDU+TAsnTq3soHcGWpRjxk0oRC7tQUV5CtkeuKKxYvu9vSf
RLicacO2/gb03gFOk8sOZHOdPJdDCt35Aal1hIlNZk+wXVehvM686hqcxCkPUpyiTqiMhxhBW0a0
WqwCEHVCXSRmWwAFsrutJ3PBP8el8TFyhi8zChI8HZ4pkQQBHw/f+OTDal3bDjTD4e97IU9Fg/tC
mr10XVKELcUMdBMIonnju720cC2WXGIuU5mHqnM2DyxqIu+fE8PJbvFQbJzaFKIgzvMzLMP+mLMR
nUPnoFPINFgBlq+6MWD081piYz+9fyiDWJVv/Xxulxx6w3dkTyUsn0j/CrDsmEAgZ3jd4BrYHLun
5+zYZkTb6WJyl1e1IQGVeZR9XpZTMXwXQJBMzMFMnz41C6rdly8XsO8qRLTb+cg2j/artZA8VRXp
XI7JqJGMgiLHcS5ebmr1u0n6bQfODxxGKflUB1fjI0Am/6aaGa3Q2zzq+O7tpcEPweNInnN4ehuJ
GyLu3ruYd3LzUOrdTJ86S/C05I0HVLV+Z+m95MWFh8Owilj3KdRvy/QaDw7/iRGfS0Mj3oxtEX/0
518+uppU0wB3tAxXlVyaNGzFP+39HPo8Iszeqx79qiMy3+7U0FkgppKy0VwoLncz1150t4aDuFk+
Hvjupz7e0ep2I6B2cMbxx1j2837RFWNPrQ5IW7Ytal2VmhYuuz+ZyVN0uiZ1MjUjYp0sDcpR4vkN
QiMm9TTz9PJ5WDc8oibBZhJdU+l8zZG5CKXrTTPszMkBoVkKcXp+RCDwSiB2/a4AJAm5FR2XszeW
hOr6XEwDemvBwfrNTWj/sigamRtQbTg3xoUvCA/TDr4IRH58P5Cpb2wUQcMLoIlQgd7zCYo6Gu6n
DhqOFtTUoA0yj6r52CCGZett9WtQCzOAFZWe5oEmeGSgqEMD4WkUpDdLSGq/XF2cYyJAPSCD8d89
oPKraeKtFkqCBKBn+UuuzYayh9c1LVY+6LErBUI9FI8ErpmVcLKrqze5xI+CnjhZVMT5JARxf8O8
TaEbY8yEYb7FxuXfc74+uu+2Z7tHPHfSg/h4C1XH/DI+zFeKA6q6iYiFUwreOfnHpC7at+cFxUk9
kl/L+JDr0Az2ryrMGbTUni7ekcGC64XmqS8rJIM7cFQepTGNYuh2vGOwpdKUvLyyXEt8n+tVuk10
qA5fkD9/8X6M054BcyvfAP/q0WfxzSPBeDsSEsPI4Te4XvXelWim3LV0I8zxmkDJnT5DO2DkB8jk
z3L9Ha0o6Fxcgv5HDDd0PQfo4SHsqHSEPYBMChH+hhnRHjtTm7GulxQPoTfhPZ23X9e1kxZOMwWv
hXZiQ/YB1m1r1edEgZr4dWtyn5HxaE1rQ3/Pp8mWK+ISNEUiQDFocWwLuaSufRiu+fQlrZ77VnDq
GDnyLXY8tL0/AA3515/5Bt/1ZNNhr5iFqjKVe0HgQGly5lQWbigXEHazr9Em8IytZms8e0PjORfO
uDhvS53Hnh/bi8japUe4SO0QnWLKqWUFG6bq3xhpZJHEFIuDC2Paxxpll43A2Y8/Yh8epjwIbeJT
UJ0Hm5fArh+/lSjVnNGaolnRkXRua2ko8qBMnqyxCdw8xtbKMJren+0RVrO72P5RqooMJ87sKf1Y
BhsaVUjUqmFQuQRCTq724o/Wq8eLFOw/5RR7TQniKuxiz5wN1FUfj0+Hq+70BrZsuGh9p/V95C2n
KHnU1e1KTXwokSgEuUUeOBooORDYfUs3YreSCbsm0uBPacxiPMmIvp/vAN9x7AIErowKGPJlBFg0
T+s/RFstu9T0G7vwzMDmwothFv9RXOGrAOHqNJmDjCblxGCBZ4vIIA9/an1TgL97HeAYU8Jgpc2F
zhD8Ync1rBkd24BwzDGf+3lUolZ2sFbKeFBoUXM/weSqkeL7Gk+t/V1PwYxYGrWkpGmOSDuotLT+
kVrWJS0L+sF0FQzWIAW/zARZnR44xaBnRURBXf3aXJz0RiC5TrGL1OuWUQI+053/AjHAd8PmoZRY
x51waWUk5+851Fql6IGbjB85j6+U29YJN3YFHixMoO1rrNwiLOXr/GuD+Pc/Qubdap+iPlGwS9f0
JeD8+11uWmP2B0vlml/Qgz55KtRjw5wQk0fRaee5l4scZ0h5GmIATI2LtS1iaK+UHb+EF9Q0EO9o
5W2mxTobnqkLzPJ0Lc4gjx4vVi5XMvYNcXUl0Xw5F4sWaqLRlnT30BKeyt/zivxSmwFil8i47HGF
jFkbwakFBQs1kGsA/8/AoY+m6lSoaK0ozIqXdpgiJAnasKXFnGFeqDJJvZHkjelXXb0f2JHNMYfD
Qa0dSKvWKUkeHksE+Bhoc1YWz7hucXT9L1RAhR/RzsN42JczkgD11crhHe7SblVT7jcXsMEf7SHp
end2YwZQ/Gk9vnsLlKpQJMIIG5q5mE11+prJfK3DGVssFbdwyOzmxVjYphDWntptVqUW9pY3Mu1+
0ctLpdd47z/kpcRCcdom7J1zmgkxI7RiVmsHxJuXCzGofKnhx++l28REDENPm8PUUKCnbOYkFVjp
+WwwhV4jiKXGyEZg+cV/f6gMkA2nXmA9zw4Gwpz2XxEzHEupZl4/a2YjrD5q16YhicHnkN1DRWn7
qZzIvKY8zCJNA0P1DmQXSWii35M8Yv8edee06sHF+wfmqT61iUzBQEy3obuKCb9QfgoowxVEKUwA
avdTgDZtLnbyX78v1rHqGrY6g7exE2VzHgN1zfXhvHiCzILi+HEe2IwK5beA826SWCIGCNTfL/Ym
R9riHWPx53zIB0Uuc61K0EdpsLAqLOWqccHAhOE6Xg5qucz+IaQuxVBIC/sqqw3j9Qai6MVzs+BR
GjpxqHaY4M+I2s452zLNe4hoQL4FbvY1VB+6JFN0y3IK2lXYF1Ly/CJ2cWYdGivnOfbzB8AfW8dh
QLSEQlsBbOU8dCbwGR382qeGydqtBlxFFlSxbPRhwejY2SHLVntTNjsowLPCJgY/B/z9JyCO2Xna
pFbE4N+jEutL/AP0CeVRYuyz+CgMNEErwR66KRd5fHmHePP5bwTBcTDUkxMgMncJ3sSVDoamEI0N
xyXYYILkPrQ1V/mOepSJ5c1OX/h8SftdiuizfSYWwwcjexsqRo7XF4LQ/E/mJ5oO6UKWodPCrNXS
AF9giQIkelY+t+CqZH7iXtvvTTp6nMkjnSygFCbT6GBiPsBcRPrMnS8exjIuzjFd0GEN3CByPzv/
OOgG8hoV/LeElA/uwbkvHB6kWerr8PBwZuS9w9syYAiixTX0YxMpjpaCKH5bapJYnFrbNaUapO/8
AK2qHQZwDExv75s2C0UmD407fHuzox1T7aSBvJZgMslZ7jYGWtsGru3n3LODe2T5mUJ0caEaa+5M
oqqTI0gELgT/7llCeB25RTP2ittltr7WxeUrXfoX2RW5jh2JKyGuIEXwJer0LChV2gbpWYmkyrP/
FvQLQXDdZLqPX2FsTHe9Pu15+FfVSZhPk2RQcUGBt8+oMm0D4V+dgrkxGUtyILwifwp89IrL+lLc
oEFxu7FBt2B3issfkWSrMby1MMAKdaPlUsrBR/voXtqlo2q2YPlR9lFCzuCThtuNj2Cm3BEj++3q
TNF/1terewKeiQrE/lupktgv5F51d1kC6Ybx6euREN0WtjrZF5RIeUj5SLaNT3IxKbfn5vu8LhT8
8kq2jYupJMmU491qPUZbjSPfGGbAw6EFxcEnyjnL/jx9IWJCStak8cm13diXqcLlq1OiajMWS9ZV
2tfnXwUvKAPGJCqhj9+j1N3YoCM3XxE+6U0DzTPk7XGYeSODxM7PPHEHr0MYvV76LBjJfco/tLCk
1dHrseKvz/pcj5KVJFN01E0jNByN4gSjIipsRSSpvfrsZvFbIgK9gk1NJ0hzJBK6UaK+t3hN+0UY
8Dx9PpRGLDDFuKWryXpbtFD1kbxT+bc0GZJQ2fk3cD8leHGVW8EJxE/B5zzLH8hLvd9+khSFQa/g
kUHNFLnF9t1pqTeSNAtBqAoyYaBquqWHkWAPslYJcGMxHBBiN59UMP0ZeRcLG+ntTr1LPjz7AKIT
Kid4YQLUcK90tln/yUhYBoQoWsAlyBNTCzXObZwuuSDoo4Y9L8nmekLkLIXd73AkQodt274qXyZx
RCsj53SWVMN4+PVbvs7bvtra8l8hOXgMgHqjpKh1+wgWE+zcD/G1ghL+asokxpLK6o1unQdWQOr6
udAX8qllndsaMcyYYumjWcHFUs22tJKy2obaH4mH/O+JbApAEL53HZpaGyEBNEoAM8MM6iLb8Nrf
OxS7fv09w/NRGzifz6tQSXEU0t1juCJ+xRY8KVneKyfQCZBTGgPoUIR2HgAUJThvBd4HIWPaequ+
hLUJo07VgmqmLuGzpuzQMdpLFO59qi+szuRmuFcOoWJQdXB6uf4tie+pjSudmuY/TRBDCkcbo3Bg
ETJYoDTJiGNX60UhqTfm5BkfPYYEBcIpXrlWx9wuerbOmQ3L8GeOhlVHIY1C+kH/Pb7u5vQWY7w+
qJkU03tYMO0lv+erKHr1aQNIkNNOnEifbikp+zG23zOYy3LyxJDU53+fFeUmxEqTMRQXNGYoeVNb
4naE6f5HbOjRYo6DhJ6KrffR5GOvm0ViBaMWdFN+ITbIj61ZrTiROJvz09ckaiYca/pn9DpPGQnF
RVOnmwGFcvsRIPLoc5Xef4D6L7GqjfWGiZP5tE75mXbl1a1wGpQOLcH44W/Yq9ESVdWR+R0HUTeH
uuPrIbsN2i47M92TicJNZTtNSz82oYvzbCwYtYmZ1dS1HOD29CffE3RJuRv1sgzwCzdZmxw6xvqa
WEkDaz+ebqvH8QITHnapXWCFf3I6AnDdwqaaueJ7vZgk+QtBV7qldmdmA30997P4Klb385YQ7jML
3iVADMziZU+VhKMQ4Lf1mnsQD6PwlqVKOocrqEWRsetSDLtvMyOAJsxDa1WOd7TT/sKf13u7p4Ev
QnJj4PHaw7fWIT6IY0qyaLX58Y+naBgRX6tiJF7YvcScMiGhIDZvYO6t2arnTUlbA4wMd16w5VTY
vc15IyHVhLvFjvdeF8y6a8ZgktjH2020UzpalA9CzoGNPJlSwY4eXKsbFpYn5hqk8JapycEygqrw
i7war8rh82Xdz4fvagmaffVXLRoDQznXCT9v4ozCRsTEnPqK7gRnONm1nCCdErCOZV4vvnoASYFK
QKQEPQKUt5WQJysLYrzNkuPXHoB+OIeelPe//KINqQFsauli4FvhP805FS7JUY6AwCgRZxcQE8k3
CfPwlqb0k1b8o5nq3P7U2Nc1GKhGufZhUdgWR6vZY/tzVnYqCF6RRKn0yZZW78ATA1FMpeNVGOdJ
uxhYqZeMKtvOf7JM/ukiA64g6qmnE0gyzsam9WJqJsfp4VsAtu5BLct5JgLwzoaR1idtD4GNug6f
oDaeT1ltB97kgjZJ0yFGzUM8wJJEggSsuIVt/qC1MeZSFeVO56F5Rr1jXmAT/9+vyXzz8GSTj9O1
mWlI0bUh1SpjadWt7Z7vFofOUMNt+ZUF+4OG7vDGYs2Tm2rMh2XpWO8h4JVJiEXx8Vf+0k/Q4GSZ
aJQbECL79ncq0OY2lW9u52ntRvOMGEiOHsMAcnqqblnqQrbgopQOdBVdnYZOt0FwnUn8OBA/R76v
LUcfkGTJayM9UirX2eBg08VS26fhIoxBbnAqkfB6SGo6cgD1Lu6qsJOMLMwhQc6t7+WNRcxwkCz4
RT1eaBSak6Lhu/HxPdXMtCDTwbnmcBFzrb0xCeE+ZSR5wsaXsC/JRkb1fE8W5BPS2XECJ4EfbO59
X2PRrHrACFY0vm8KSC91+PtCk3tnnpD1y5ZzNZlbdcNm25UmKrCLOlomlu1y2SIgmDJL6/20lbxs
5TFKDqYbWTbOCqTNjQhOb21jk3Al9NmAYgIYickjy733/8C+MIS9lHwP6BF10iAnKIZMA9PzYF+q
dDrRCXnuOlVTTk+uqXJUmKAsKfI/nIN2A/6+MV5yTD6j3XyhUCQ+dyzkAOZng9q8L2XQNh4SLUWo
hSLeElPNZ6J18O6oykYmiQc+gcb1ZCQX0SdtzbCSdwvHKh8YHDAw54M4sxR0EEsgma1laQXAN2+9
dydUbBbpFMSn9QxNYAcFPI/6k5uLMWUQWodp3lR7xXuHqRNtTYQLgknbe0eGCSuT/Zkd6mU+D505
aRLdFu1TlmvtqT5CYbhzCor5c3QHBhvIk2c1gXjzVQHKfDYrV5Xpu6fbgzfGhVzZAqhpkGNhdMn6
V++oVv4tRAHzhsUApK1Ia53uf3lsxhzKbNIjUqm930M+xlYl2cEKqATxrwRwB4TCvjrq/+3m+YK7
Mg32m+Q2hLQ2T4Hq/aY0HvvIAINBTGphKYQe6YEbPMRdl1vtkhqzgbzQIf//mxEctGmVGjWLl0wo
MfoJCPZ30Gqigz7sS1xDcXNhXTt3fkOq9AzTaP0MuQfjG1i2u9Zt+uOwWZpeLFBxYX2bn4DDDDUf
7u9l/ScQRWGPlYaGgWNeH5dQH65DUAZIxw2mdHFCENnozb8x0S94mO0p9V3ZAclHFC/QY6eX+5eG
GSeQhjra8aRMCJL6UPYxqy8E4tNiW1rUDtEVvopw0jkzyO+1h6TH0uTy0Tp4s02aSLGaOgSXjG/h
/Y3jURIPYt1ZCeKoHD8HYFaGKAnMUCGAjR7VW3ylTDi41dMXwRgPUD/uJDycc4ZJQOM1R6tgNklD
/B1qeJYmioIAX4Z9gTNZzEohbKuWd/V6Q3HhSyZrogDYoeYx+jRhiEdNnoLJehWkZI2Um518/so5
bvBvjwBHFfF54h3Jt859/4JDy7UWgaxAm+3choAZ4WrTzJFpPlnrFygqYUCq0KNhIYHbp/5H+8J7
E27Qq9k+/Bffra1o0SDPiA9R6rXmf4NKwh0hbOvCDqvZ8z+FoiZnLuWJerDkzqCEms9p4/VvnpUq
wQCxZs9ug/swhVsbSPzZ1FtQULLZJFKHduKSkZemg7WDBDVdmOfwcpKyjyfmQxaxpAIYKQf6U8JJ
UNYkeTOtFJLHJxSwiAsTY36Vpv0yFLN3L7thPBWXOuTvWjbMPznx6xD2xu/MmKhdM/c3T99Xohqu
PMOCZfWYlafHg6zMU1J13MeRJj+POYDgxpAAuI3syXwrJh/5R7e28zIwiDQNjNB+b37r3OfABBvS
tnrBSPWGIx3+4GFRwN9XbmN+3eRKHaqyaF3viBCmv0UIDK1txoRJRac8IeHlk31Xrro+E6nTvQTi
dRF9cgIxSFhyQGyJSgKRVi4VtBWoxaT7C+YffGudWdWpvgiqrI/ovCeTGgWNb3cMvVg1lS9+oinP
4SpvLWEda14fTBeGu3Py8nKT53ZJwWUWYNDWxMveSVfQ9t71n9SjhjxFlR3htfHUkI4H1k7sF3VJ
UrRpZSCVS+qnzCrzathwWMxq8YohTqfgFr0FvkadxXjccidjAmOa8fa1y1AS1Mf8dvamJoUApryd
Ak+jGDfdOllG+iPRLmHxEFaioLgXK+HA6b21ZlCycP6lJvOQyI2fMlvOq8k4GdV9i99UXEx1G0u0
LfSBySkaPgIJWDbkOa4bzcWM07mvpQz+HaNkLSL7Mtj83iYMxZJZxWKX27dKER9cPNNho+rb1t9y
WsukjP2Vpvm51Ng5pSSUb9iduCFVHAqAsLqaknmKP1xvgIm46S1/Kbn5BGKRxixzlMi/9MlgXlyd
FXe/F3ULEyi6t+EtYg3iiNxnt3Yjo3UZH5xN8WP6LMkJI08EFuKZIixJB/RQDfXVryaXi94WxBPy
U5/i+hmn5JFTJYCqnNSiJAul2Q3v4G2EqTXq86tAnA3np4sDKwY0QajQZNDdUdgnOZD/dJKpiNNb
5GpyD1ziQMhAftam4PCCvE+MtGiXwMCXnuml/1AOR5yzaF6Q9o83HeD50tu5woWdFKWHngdcL8q6
1NAAoLKb+5B3e0XLxG7g0JDa7YPvftiLKbBu2qwf9DOuqDMocrYiX1/klNDOz2i+9/J7gZ47/2PJ
50+zOQWS6R76am0VQcGru/pRF/WxHer5NE21hfKA6mbYpwQ+6gqYrleFTdfi5eObccpI9gYiLc6B
9ej674gYTjVApqb1zGtMZ0CtLoK8mVW/sjiKs5pMPXOGM43E2XOgFXFWMrcqGx5PRZ6zZKEbmbzZ
tDtp32mQ7VEusGKmE1JWKycAIkx9w+tnp9PFR9lAlM1zHzgyiyQDDZUvIKLAWR09s4OHRRoqt1/e
xhSw3jWy5AVwamDBWsZd72I8nHA3nnW8WuaysTLmH+gPgIeEpgE4XuZalnZ6mZFKK+7KEmvarSup
3yaykDLFR+nftCYrvpGmqpoI0lGC2H2K0bkUOGHh6zNmwCMRDpTxR8nDd881hSe7JEyd5Fx/Gp/H
sTlUKoJPBT2O6gd4NhE1HlydpCO/gi8IElY+AqnXnLlVSY2apBK+cmuH0BLZVLEQUK/sjKO6uVVu
xiCphxtz54vSsWXrWxmd1iNkr8uTcYpb6qmCFsYkMYdw83X5eragTPxfFCvxQFKTaDN59Lktresr
iVDbBsM57qKvfSHDMPmTsf/YBQus5cium1MV1/wzzZGOe2Z24K/ToYb5rKeylw89XJb4A018Vdb0
OaPADFX/kFrlsEVdlMQnERjUibRE5XO+5FoRJgJdH1GtqGREQipUgpbZJvzXLRKIU3+K7W3HNi+Y
0w0RjxxCD4BqBqyM3LnVtUEyxniTQbvIAM644qW0saI1HPJQJBQWL/+OPrsoK5dOeqJBmjhaT3C8
/jkLl3ZRTxco9mh4Q9dCiLTfC07Yw/GtRL0ipSff2Yo2IPKFJWq5667Qnaj6lRvLdqpJEEpaDdEX
HlpC6S3MoBqseeqdFqHOgC1rd6+4DVLXdiWDuGw9o9y6E4x9hkMGWdj34khjYpVANcYmpG7gazge
2MFIqHweWtxHW+3GKJzMrJBALHpVoqS3MyE66YG8Kg9I9xPYoEEFZq3T00ZvN2xNeM/TIIck+XSH
9Yu6XG8Rg3W+TUT0m3CIIjbEjL3NQem5lB9btFE/1I+af4WZtyD6aKbGIMfwyD7WObHoD/cI4S4g
D5cLPv2vg8uZMfTnaH9rQGShT53XhvnDXl8Ara7z2sEHluNffzA9NkQD/VQzF873zS8NuGOEJhwn
SVBn61Id1fxA5vn/LdMlH8N7x68opYBKTtMo1IsZe4UYl2V1ldO0Iz6bhLMYzuMLOFbP4MuBSFlU
qam+YHYN/wpD0s/WcHyb1jHV8qhC6NDYdBEgIYZL3SG6zRyKvYbJviHMBeDJs/su5YF4XJF/Y0qB
gm/NUtUOeejDqKLSgVFN4R+jmaLNXJq3JRPNJnMg5Srm4k7IsuVOmKczkAfPk+M8cOOJfo69gw/m
e2GyhmxOaXISlbzbGafLvT72DRkjuMGjRqU32Y33tgM6UEFL57Vsi6BlGtrNc2JdgvCGvsEdhE6O
d2BxCVCyuPAyCzbcDrVlU/DMf+BuZ+xoQ5tmkTl3VZ4Q4m9OSkGm6SQqMqqMUh7qTMEmeUtdYQ+q
0DXXIUG3z3euryLwNAu/sshOyJ/CuhNrgJI1Y4k0mG968NEyN5avsjDmjYMZqeKA12rNO8U7hqW0
Cv9tvRY3bkBoudqTXZ8R/mDSCRUcb29k0dNuJFLky1x2KqOKptwnooaJMbS/+2QQSkdXzDm6yC55
soeVN9W+ldYRveNrvFy9nW1L+kz/go3unCjj0IDrOhCPF8iRBRk4kUFo2u3jFx4sxFc9g4VoAUbv
7zHQz5RFpquSaMxO4wPWurVFz+0F9DP7rFUwXH1LrUakLpNO2OcvXFvPufFIVw/eoNR3hSOlL71m
ZgHGybKy+m7hNPk9EjvAY4MRKaUo7vt35/gaJCQNIf1eMsZn7knPIZdhw76DZ7cOTlfwDAPKCUJ1
b5rtL8Ptpo4/min6ftwT2du5cOe9O1NdS979QexJIGD7rEGrb6j/56WqSLy8FljAMABfaeTmSxDw
63OOD2npRRxkCymESUIXmvrUEbHWKZFxueR1RtgNVUlaDo5X9f3jpIN4RgcwKU9dxc5Oxs2vhaI4
0FBBzyZTCzu6Ke/koEMEXSYVvBPm0V2WIwFxD9Yp/vSnfwPr4ZBWKSsQ78rJCxWp/XQmwIMkkbS+
J5N6n1cJf0QTZRFh5ztoOTV3jjZNJaFLTrQQtg/0wzAiqcnokwTiJnKG+6dn/1hwR3lgm9mE0FuQ
yDGK35ibGgE7I5cZ5ZKN2tw8drFIy1kmkKzGpoqd1qhsHKT551+R8E+sDWez3CyHhdqpfWfrppr+
0amoA/UQihOXf0145kwSF8Qy2jMR+V1MKStpExrEPUVwom79LT0Jjp0orH4PSFQrWH6aceyZT2yh
J78yLYLuVnXDnsO922ODzjK+9vWwtscPNVFBECiwtDBB8J54/kzMPyd2RIrzt5UN8h5BicomhnpM
3j7aaYfBsdNbiEJW4c8kIXWS0UV5pH/TzPgCqXHp0pZxI7+6eCeac4th29aK/zOmGr2c+cBIdSnk
TmgA0TRnIAbZ0kOLnW7/P4vn/HnbB6XnMPZU7JfUWlzb1Pl1wp2KxkUVqofS9utSDc4QudYaLrJN
v4YIHCJevAktqqfzj49M6F0BuUKme1ZycWOun0zZ2f+aqLIIgjgnkkAASWFC2i8C7IZxiPU1ZPa6
yjrwxRONlhmTV3AC/NsfT8ECglRyXi9sJqTPBfiYfuT0GFffFlQQC3TtaQYGWORFo2qzW+TbdnLJ
D+3aQLjs4mrgkmikFWRXz25hPZu2z6Zng46f3Nv+0vPdC+TgQoaqiHEy7EkupimqwjsnB/g985jB
Frr5XhPls04ySSbb+xiDzSu5cyNZNUd+sHdFs0tZyCS8esN/226OJ3ge0DnmGnHGJ9dAWJq15p9P
KPE564o+PTlasJqFVDXkJH6Nn3vkCnl07GZF9+ixS3sbrU3AiiEhng04KdPUJREnJ7ovYWmgjXS7
OyTQGDo/cm9BuW2s5gAlVmf+eIHBY0tX/WChyYptADSskf0nM4BhNBcKPC9j5wlJB03xkvsu9PQw
Dn6tMmMvUxkpB7QpWmDcrbNNNSYzbDm3UneQ3S22ujD/1i+r1ZD+dP3Rag3fmqnq+1GrbeQXg9yi
B8W8XHGjl5DCdTyaXbQ/H+wrVdScnZGHoFEk3ip5ZX6WSj3tq3w/Jkel2mW5k+aTyj7m5bFCfpmx
LGd0VNzCuvRilGUeEuzXUglL2owAdfapZhLlc5FMT0f0lVozVXl9NIwgN4rBcx5ERoSK3m/1z5tv
xk8rYx594aJwT6Mu5kq+wLB/ubo1w7wSOSH4qYUr/iA1KrG/WlMaNjJJxXew3CSXkGug/gt8DI11
O53Dr/MF5x9FhhuflMQ12uIJiuF6bm9iWVxf+A8fQ0uwS1uT+mOBd01UtPCYdS9ZgmvAHUwnbxvU
QEzYu3s8Ios0mOir163aKRAQ9pUwiVgqgYrA7RWh+pvpqbu8LyOzG62/lFJnpjBkKja9Ons7ZT7g
HiSHI7Fgouz2X8ZOPKPeD1tX6ZaewQkSStdAUpatIOHsvOublrrxPy2p8J+5ErQQRBHxmo9p6qeo
s9jIwM94a8dEWRFJIJv6VqhMpNTAnNlHeoUcER8QI7hADmigSUB/LueexmFB2c45Ds6n8txTtOHK
U8pT61TsjbcxKHL8+HzdYxH6MHrZkRJivBkcTZS209EvOOWHAPMapi+9z8NQUYzEQYC23NsdX+yB
i15pmbCBwrm5XeIhFhn2YGtAxUETsCJZLwJoWQPn7YB75gG0V8I0lBF3xsnUR0i/3PFhGs0PpBZn
QfGAWzw9LIlmhpOmeMK3ULzS8eStfCrL8ZDVNeRpTf0WzD5O8fqeAgvsubjilRb+bP7Upu/ipBmG
t9B3Y5NzlQMrHWLkxb22uhTKp+PoEtHRMv6dctHE2WjdzYX20cl0QeblbGtkcbB3B3125k0gmKnF
/PVbt/MQhT/vzeYHZ9Mc+PkKfc66jdJychE8nrMT3ex7p0QsFvyJVE5xUT5hm/N5GDEgC96kVBo+
8hMHgB0KEZNdXkP+uqRNxzEcRIyiNL4ZM2IM0MJ99cI4M8b2WL/mFU+geeWLLZu1E3JK5LzWx3rC
4+DXlHwwGGUR/GZwPvRPHcxAtUqq1ruoq+A0CxKK971XUAI/CH24TkNuMGgTmT1oHzoccyDwkNL5
F2jI3z1vcO3YteH0uwXyA0w6Fy8kOazAJO+PJBOIUivANddlHvd92m/hUvTBzWW0a6DKximmDP1c
I4suVzFPnZIDMSvn+vaj8NijPttKXiyPzWKEme9ISaxdEi405ygGXDbYVhihIhTb7ep9J8GRT71y
BQuvawB3Se0P2x1SNGKAW0c/6RsJJerJEDpImKWgZWdaGR+ZKi6WNUaqQUCsfyIrUVy4Hbq6PQlQ
iWTKZ+GagYYzF5hoA4E5PIKkX6YiUncbYdTnNChMTg2ZcbidbXpdb9F6+ghbxkMsAkICn8vXfCD/
A8O6sfPHtPj91i5Ab9f5lVScArDpWLTl7RuG9SMQUvgR6VHFStFz3qmwLlosJG9HzEzNmAV8tK8I
kBnPFwrPAclqrSUJ8oauXRmzC0vpDp6zhxnNVMD19Apeikr7Q3NK7RPE4h15mIQNdwi7szGiVjBA
zxu6YkPVCyodfIhdRvUI0OX+VTiTOuTWyqtiYSvayqoO48XR1cCTieClrkd4xZ/HU35sbNzOh/6G
59cwp5vsRZ4+ILAaqEbe3/ilAgilLKJa5PF0EGWh2wxgjTqkrYSGjKsnuEyUFKSgSIuwBEWHA+x6
9AikoVqRhPxidP2Q4aFZ4sCuYHJ2aBLiLlAnitd80ouZdhzx3itBtBfoCrAKCknRybmKKj9UDVMe
S2of3Nul3s7IBFA8QtIcrfMLOh2e3B4uvuPKXeeJtZYYnFVyc0q/W906Rp2znJjhR7LdHf0fLdND
mfZHT5Hpg6uR6eowXVtjpD8qkPKu4obgnjqjN9Yi8cJfDph/H+oRTXjCHgf9q1/gASMoIHEkexDd
cT8PqJqibAWN2MHLM6anfTuKTdVkDHjm1bb8wQH/m9E3fB5U0qOlmsmM4Fi4f/GuWIbLuHvqu6DB
XTNHKtgcvsd+dv6jeEF8iontWny/hb7TGazQJp22/z6pkdr4O9hiaXYuZKg5aglOpuP8hoAa5gIs
1hdqcVWrn7dSvp1BZjbDqzaNmLeKUpPuJSS7M7Wr/DmSrAb/83+5ykaRLEmdImwySNtqAuTfwOiB
VHXo2dO1A5YzPAcoHoFuS0cbjf8O7BJm8ZhF//tTsE+mRYVFmTPO8ST7rj8tF4pFzti4XLf/iThE
Zib3c4qYyONgODMisoZt5ipxykN2IBRXBl/4tcTIVsdxa0UcxvPwjazLVZ62y+U5x3zhcBfweLh5
VidQK4Gbv5jTyzuEbVlcxLg6Kwp2ZonORlq6tZFUFXbUUpSmpk2pbPSeU7q+00x/ITL4rDxcijne
NzFyMoLuGn2XcJBca599jwXi9+GjiHn6icdUKlHQ1Qz5piBgiK+rgfo+NUT/pvd454lG9ZLXsHlD
hYn+JkmDzhxQCpGeZVVuii4uhcQ/X+X9d1npRo9tbYR4VA7nEiIXL6cZYIqshc9r0YHa3pNnt0FT
nnVc8smDBEml439gbjkLmEcLEFnv+YNks4MDmUUoJsZlAYOxmyWrlYK4oTyKeQWwM/momJBx6KCq
CSlseuwoEJ2Y0E+OyZFUpj/BLwBh53lKFT00Vx80D5VqoABQrTCnmcERc8AV/xgoD64LBENYbDTC
3WnEYVkMZ1MoHQZcsp0pXIjc2owCsoySYCBqX63EiMuaAbebi+46BIB643qvDZgULr1nLn/B5k9r
ampvyiQXMgxuEe4X2uzwQPiCf/t5XhThjUtyB1pTF4GmMfPAwZjQB/5LYq+tnrzqyj7YHyJz34ty
tESNxEHHfOYnh8I+7jvIhQ+2kwxQtAeD0p6vQKQZJs/ULLIYJVddFg8gxfKBRV8YEMSVvSaVloWH
r8IIR9/P6ift/W/gnvNJQIh+ldtLIePGU7FeVokc0yoE5u47XEpXHZSQhwvhCNoGIVcPOGIuTBo9
OcPTbuOUuxnsokWbdOtD7oWycTD17ArsKf5ZKUDqG3+/UrkvTgXUeTu60DBfOdlPieJzeLJyFma6
dy4J/8myt+LeYQrxNGKjqkJcR7fomkNOUbTnT97BhgyJNEQ4QavMy4g2YNGKUq57wx+QCGtRUc6z
1oTWbLaOiJbEn/o8K4ojH7e3O8LAvtZEndyxs2N3FiJQQB9qK38VI9kSo+jCbK3mDIHapdENyhzi
tSPJ9FcmvMXoS1dvi6vrN2P4IMu41Fh5epV5TZTg5np/muyuZD75lv8+o4fwQFy483F8o0P2mhAV
KefQvX2BiqxsssXNHzviamtyQEFiLW84E+1L4mxo4hbQa8cUGld8A5elL+/8ROFCtvuFp36R80JU
mqmUR32EerMaAtu3Nbd4Im/OCcmJFItWjJwheQwVOaydNkg/YGuEgs4XWH4A/zgOkHX00h3D8wOG
c1vH7hSqReyrinSeIakwce1RpKUGR6RoKM0roK38nqFH/ael99Cjes51kS7HJzUN3xJXzGUGcL1f
gBN4v/k2BcZaP0vZ7e42CtR0fDDWoIVFcl9GSG/m1g+VuAkYmIpEWAzlUtxktQ89yTGdxwlydR8D
pZPwxhEXtbsVfXswTDdTaFdQTWcDbUveXUJFblZc6BQfh5er0Zr9y3FuzOKWSptyHW5hwHpMrTCd
CZsTP/7p7YR9xvte1z2VFqtdHOvMG0NH5GhovuxhifoOsW11uTQl1Nmu2SWtjzWd8CHM5CA7W7YP
5P6LbkGok6EmHgrrbeErbL6PAVRpgWk+Z0v+LFzPRC0OJC0xCh4tKgf6wdXBYJ380LGTbhELqgbE
bizlgdyFxzhLka/sOSn7LOHqmyprYoqTtcREu7bx/VwDDgl3jMm4xpurc0OPmRl65QmCHYkFcmnW
mUbKhSbGLFgE83bvP4GsdTnVp9hFtRZrbNeviXttHh2BjCKbSQLgeaPoYgbSNEVoq12ZE4TAR62t
Qf75sQkVLFwcA31TdUmNBWehp8tGI5BmXQVlmsKNeIbP46EnGaQZ8tRWCbuhFEQZX+9BQK/G3tLm
IH0aOZwnAbUQOvjIHB6USxPWKEEsWS5CRLylX4Msp6IDQX6qodJNHw2SaTCskZ10lwdpnB98gmVB
ZdkfsoBTkumTXSEeWTeopCxIGcYShbtrdLlmyh9yJxT219sLB3kU7MIOydJTRwjRWiQYmSy9E7VM
GWb3kOuYP1+JO96DnlBvbmoVZAn3jAtPhY5RAwjNkPMjCw0eEsmKg/NJ8YARkhaDhsuZk15fknjz
yEhMd43NtkL499Ut1bajuIzyYcrhJbT5hFfLFK3OK/gwkmtC52CxExrgCCMoc82H/VErCIn5x/pt
15YfzBECOtw/6/uVO1d0b+o+hoGTfXjlWND1DEla8GlMnejoFcLNq3MqSfjL3iapvdbhljd3vyp5
VWf0INb8xPGJOLXxzAIGVaytYa7hB0n2Y+wl+9TfOCZfOvpqjZipGzTWLY8JDAxMJUJn6qPoXxJ2
Lx/Aru/mKK0SMkbeNUCJqz3fN6Ofwk2bnvgoVMIKsRGtxeGgGP9GZ7XI63urKjPG8arNHM+Vuykh
KgpGoQpmzigO4DZpgDSPOOPVWvY/YLilENhPvheN7HHdzkYZ5AejNfKNCAr9zXDfeCp6m32eJ7o0
Cxg6dFSafZOPHgS91ywAcsmToS2gLZryiMU/FpFXorAe+ULNwsuMcH0uFdPSmf9AbdXhtQ/JWhDr
ER3w4KXcwT54faf22LpYHKECAMR6cMlrzpAjcej46jDf3OXekcxPI2eItYD7rAgdVypdDPwaf6gj
1VnACk5JppMTEJHTSiFJTkFkHbuK1S2mYBvt6U/ypA+l/mG0uAIplN9/6XgYNqXWtThWV4sDN+uw
tXsb3li4NIQE4+VpmBa+BEA06hOHvxV/2A8uiY58J2NomfdpoAi3TezE88CGN/3GW4/9nIiMosk6
jUzT0iv3SxC/Y5DZpZ1xC17ohVB2Xdxz5t3sjbVgUvh2tk+QjurLQ5xFmkBCS8SSaBIAYWG62vDZ
C2xP9SH3o/m1e57ka3M1kXK+kZKQsgvBkbfMqxhkGoGzRXDgBm965GTT60zHo4y/S1hw0krC9QZA
Smh/DZezdYeuvlUduX6CDa8RWHcaHR459aGzpXFdTQGT+9cVASoAI/oBSNwkQOhaXXdFcC/wwtLJ
iC8lajzXAW9XlaKdayp6bEBOAeQSXXq4jGwm5tt0TcCdLPb3ZL9pWunPtpAIWe+KK5pd0Z4ToBJX
kQWx8885U5lnOXmCD6svlahv8Q7vaiQHF8m/EDmqaO8cj5MTxUz3fm0+3ZGG2t9f6yM7xo4xCpWG
ecbb2413xtRiLqMTyWMHCpRb6OD9zJDjOm7eegY2K26mw3m5KspBMjYrc4mp9Q+apxoM5aoQxBfU
hH8p/ePc7cAxCMLblBfHi2XAJXT8jTPCnZZx4lGxMBDlyRQcCsgnPOsuaKMBJKABTbuEEIeRX0zv
u81mu9vMe6xrfPJ/Yg469OEwKIhcJvGlqwl/v/fpvTqU2zUayZH+N+VTGUfSZvrstgAnzcW3eUw8
CimdETTE9eZ5NUXoZHBwlxI3wcl4TPLMyVUjxT5dgNmkZt2xJukM+K8mnUpFzEruXIRvKvmKj5nW
/PTlyHVKffwC23YYEuusGAyCmbaPGWq9nJ1j9qkXfWjhOqxKJRHvWB5nWeuxw1gHZCnXd/+Um+yi
sb6qgviS7Fnu2aQ2I5M45mSUpdgP949NIjxuzcqQg+m2TdmBsZ2lAKPeDFceK0hgl5QE0ZP/rw4M
cGkn+WWwF7UbuGvYOWL2ReocNYekIO1MQVuCjGwhrRflb9FAqANHPdpNZucRo3wONcqmW++ktdE+
pLC4y6VDsBvOU+i6Dni7tAQbzrY2U5Xf6scP/ZdQNuqP2ObcA9I7hu5TTzSjTwD+jS+Tc+/HFZSK
Qqdn/7VoazbvhoCKlRJ3H5RA5OfzX2GXjjnvH8D381cLCyjfeZhn2GdxybuDGGnV/ipyybvjAPjA
sCWB4/wlRXcBOIm/hCfvwp8WDhkpfHIGgHMyGRUeBSwINYy5NckXqi2WevnMYiW7IpEsCs0oaIyH
XBzDZvyvLm0Ul0PjDsjDSSavqhd1VlJekFQCY8ffFb78QNMZvb/BfWiDIaEZRX88Sq30LWXl3yUg
6/rC/daZCWSaNlUAYXj/k1LtdOHmCqspPyfKVicnfnF9bGu44zYfOq9hZ57PNAOkHUdnbxv5fwR+
mwJ+XuMD9JQdU+vWxz8ZUcJateYqWHEjbElpo+NVJwRBUcP6Y/U71sl8ahICk4laXZ/lbmUlaD1h
NC9a5qXSKaLb94+1rGrcbrBROO6u74tN1CJ3NOYBcpp8gL1JuqrKvFR7f4RmAUWIr5PiM6TmrRgb
KW95oCmmQcFz4Kva2iSZPqw1hN1o+qnwBO1MR3gmL6nAgPxKUw50pxSpGAe7mP9I51ZKaULAMGLT
Wk5/ixAqW4MsyYPOgc6ViV96pWLM1W+130D/3ozJg7hnNDZTaoPIX4KXaIDZQFtlHA50w8UoTKK0
VphX0ZGT4GzrK+Q4aigGoR4mbVryUaq+lvIOn74RqsX6GVWDXClNk8j7XGAqzLD6SzSM3oGYZ79B
AgujQnQ7OVbR8poyiG6Dp2TkiTRc9qnWy9QPczmJGOW7NCtYPVWjygQNZZSQSHtEMCaG1mXxm0xg
XeL5XteeMfPlq/bcMd4vwVa/xR+/3Ink673BeuIKsJF+ilwNcM6bmvesR6d8z3se572ssJ76Fn3v
8SBO5yh2KhDUcnS4zQUlzjX7BvOYObi2HFaZ+4Ld+VRAxDN4u/fT/FZLL8TbN+/qM8VgwfRSd6/9
UCkGWp1Ehdpr5RbjW6N6z/6+h6N+miyuNNG/SG1iyrpLkE92tDnGl6yCKpk20P6pCzvEhZEthKFb
xuTvBl48XKCGIClLloLKaBnvejcQOGyihER6tCeWP5P8Gs1RpMIfFA/1w3uv7qCT88lQ6Q1HLCbV
3/eXFYFhSM0wFc0mnWtf0OMZrKxFikI2ee3qNwGIuAUjEJTqg6UHcN5Xt86jbhbAZPdr+cl1GK4l
MaE+Hb9SFryWNUyuCy6H3mO78vGoAhRx7g9CRTX3+G06CEzVZk3e1TZmjbKaXPhDLSZou+Bkhn2r
j+w7P/sL4DGVlWZcB/SukXdjxqQALu1Fm9/dnb5Xl54hxtZJ5a0Vz+MeDtOGw6DnTyL/Sz8a8Bz9
s6eZQXbfZnl16tUMAbLssmSra1Rb+9YucwpBWP2ij6CIDLy7H7WBAwmMsmZO4O12bTvoORyKTWir
6ocWsTgDh5T8XsWt/mNC77Q0c79DdY7qiEnOkrTQsEleYnH0C3hmJLql+xkuwjKFG8XvUb3ypNlX
Mu2DFWfJ9KaIF3DnZielB5xMyRBJZNbroO+OptqLTaDEmS++vmU1xym8sGEIxGI52gi73mOEEFMt
IZ9CvNvQbfFb0N6w2cd21RQ/NCTjvawZgasFj79P0+75Mr/8zc0lY1QTnIySWgFGl73TEHS12aHz
ASX0m/NB6cX9WjjRJEk4jBvncnNHb70q5WvQXFafaJDqAVViSZ0D9A3HzBfjAa9P1mysb6ABU3GB
mWuhltnQQYdGOVoG0lRNKkVBBfY7bN4M0t8/asJTgMGsBZbqb1Ndu3PexsXwuWjU7sKNtB4AjdPp
cwQy8+46RPPQov67+Vtj6+3NrQjlTxYDdFEiBR38iB0oJzzZ/iRi544SexEpESguJhqszd/21GS+
i0dmpyl9zGLPXgDtOg7Cs5zpmtt1Vi/4uI+gmnYh9bF4PSd+V908XB7S8MWHCGB+Z0B2LsXoly/R
AJnS9NWiUEEy8l/NapA2TszINhwNHZ/R/nuS2r0iFQfyXK9G1ahVb0NQr3YwB2gyJTNDYNVWjLHu
22Q/quW8tyR6EjdcfA47i3nTF0ltJlTt8DIlV2JJhR2nDaLhFw6RgA0njZrKrjT+wwei/7BfRlMo
Sr6LxU04N68UQ3u4hU2Zr2RuL6ilQwWbb3I3VHtwERp2iJ9Ok/ojvg+12aU2vkUSGnrsyrsn2slw
FNM2PXQ9WjiAr1dGn4+uczPe0VGEnxEs/bTTho+wLDpRjsAM0KXr+CE9FM2aDw6z3ezZyo/VnUeQ
6JZqgwWMf/Sr1Qq2dLUMRTEYgFR9kLwBXot1FrBwMe2I5oWgf4i02vPd3def18i4ovOJOKpqsYsk
95/VYcaUfJCup45SrP5DbuPhVrsaD1OCBvNgC5j9L/DrFr8avP/tBMO70gRqU47NpBDSjzpbVl/5
ty6i8mijQ3qr+2QnELpAKzF1m3g4fPzr46wQSTv4QchAv1p8it5d1aTGvRegNyIv+DBByAzzC/95
tF+dmgEm8wZSJZnIR/pi51ekfjMxTxDKVKFWLlQPlUzIGWzmmM1HX4T+hETxDa3TqWgAsivsfrVI
lccL66Tv3AL+QmRoR+mzr9swAg9wYK1JG4U9r6xP6VhIN9ZhJsvIA7iil9pvR4411Mq73ibZ6rqI
TPGYCxZQIyd/Z67VN49DDvqGcWNmIw3oF1xr0i6RU7EVpiExzW3QJO1JcLnZHBjNPfCUWROQn0qU
nYRTkEFhBP4DHoih2vpT0OkVeV9cr+jdWYKV4SmQ44+DLpBuFv7YcErqxzJUlRjMc6p0+wBxABSa
XR0xZvFZrXjT4XvoxzcKsSPM0FyTpuO5uPPu23aJvzvJIcDqndL9pc9+biZSDDDXMo9tB91Iy1rD
D9FGNztqzMkB9tN26+VLUWLTH1X4riTqOdabWpQ2aU8/xDpT3fWYg/ZzPjd7jGP/VlqwA+icO2+V
ORq2VXcCqb89ylELwCsAHxSiroUc8KY+0sXotiFfPnevP0POOHSUpv9kcy0qX2Q4Oz13Jh2+UQd7
CjUV2Qbo6qY5te6XXBGO8Io/KAelzNUurcwaUi8NfoDIXyv3Iw7cCPid7Gru0S5EFTicZkg+M9h6
Yi40N5pcTAevm/TbIz+/qdjneRuqfm2sdcVSo6VQtfvOzS3vHiWiBOREN2NZMAfg+0/LIOe9+FeX
81Ift3Xf68D1ugrYVdcrCovnoa/ga97LFqfGaLG6s//HCAnHDSbWWYw5bujruSIuLshee6VXpMKu
dJcTAt2AWrOXjbLNUlKThWIQncDK1t82jKVvQpTbd8jS0zzBLlcTUj5ITocDAY+MSYy+SmMaR1fI
/yJYTBsfwivGqG4Xq55zEaF7yYUgXMcFcTNXeKyyK8runEN920YIPoaxlb1Xm0kXFfDzXeP3z1hu
TGZ1DWjJ2HhfRNpT/nuEdS5ZRIFguI5xAWe0mEEl8kPtz09OG6pjbictl921gZFmjFStGAV09Tpd
qytxn9+yNkm8eZ4+dwTzlRE22c9FXuzDf8anPbWD/u4KNNofwscbzRFQI+KtlhRhw5E+Z3LGKB47
v97G1DHqMS/vFy8BLOyfQaIZzgvW6jPddM14/knM4ouDFxuLXsVABmCnGvjQEXDwf4fEIjYUWEZb
T8DQhTFDTVeazRLWba7sbgprAUJKkcqnKGGX9Sb5XvG675ZTjklg5iN3kR5zNkZGB8Qx0XmT0LOv
rXETCHjgp502rKxoWxnekkYtGJ6Ta3x6kL2YVcGRZIikc9CXIlIgsqm0hzvWO5X+rf3eD3vIQlWu
8LNVnsCE2hKLgbWR3EL0oMk1DPUXtQ8SICBJlXIMX2srne1YTCLrgys3jYJCBJlIfSg6p+FLzjrK
mu53JkjhoXZMsS40jB3bRYH66Oj4axJb5wVt9zG3NKqm+u7mb+xc4PLDfbJkQCRFoMOjUYht5VqU
kSvQmiHP/1cS7hDLn1yagRmeJX1W5BD+PQ7F2l8NQx9LLF7oi9Nh1JVL4QB+fBCLmWVVy2h2Ph6G
8b0nF2FfCd/5+ourS3nSRCKlrR6ziRK4wVWEjLtRt4mDynSE55m1STVLIJCVRl6R4xpqCOhjVsHA
RA4ntpEvw9tXrizL3jqwebClCcfchv9TdIp7z42NmlPcXdncsN6llrh3URJCg/NHvgR1WgTXnjUn
bnM51v/ESs7D/82R5v5pFYQrbwI5X8xhRt7Xx1FjF4jl+7t1/dgrkaCxYsl6Jog929emu8xuwNIo
GilQtWsFaCZ0LHpNF7HAtCJEg8UAjkc+BvPdinoLkiy2269Hj3v4O4z+aIx/EZ6ye0G+Twu/Nq80
ynATQldV2yFPB0zoPDOCiUDClyfT5tnygfKoShFWerQ/7UD+XsbwttheAvIiVCvcNZTj/mZsVkmE
puRcZc/jfsGcLqE6hhPtocv2Z5VshTGg+9ZZPDPiKij/TDznAk8zC4UruPMDYj5SYw4grRpYYwNJ
PuDyQ92LVLx6jItU3456/0sNxxhxgm0u6EWyDsehkdF62waRi/Ioo+e1fqKC/EEdp+swL9r14Fir
7P59uy8UDSYyChUiywuTBMAQHw6bLLqY9CwZAx3uI4VcZQ5M4+x2Ss9/ulq71Rz90KZEAG/Wr0wf
3yC31vmaNdSDc+abg8tT29J5JSTwizgYTeFM6C6Zb7DQH6zoZc5CUhBsvw5v0gzefz8utP3cF72f
nTA5YJVWDzJ89cObFwP6iHoxcVv+YKZcD9RGM19X5sdESQ7ww81GhlG5me/PeWiEg7QJSSielgU+
7+jblzOBiEd7L1i9G5Q5Zsv8E+xbs/QhbG0paEjo7PlCsavhKYWFjzv0HZ0as8FwrDt+iKIyPYHl
Km4VEvhqKC0MxFAgHO3wnFN2qcYjRCmqOoPKCAxbLkdbDIMwj292P5C7hb+2h3haOzguROPmZ/5v
kWrPm6NsK8NqaK2U4YJYyai2Ov/O7JiE+/zAr4TrPML1aGZ3LP8uLIny5BNB489O7DeiwHLSKHQM
wmoiIcvFkKlCMLP7oGgbZHfU7FIlRi/v0rjYFQdaRknLvnbHcc5tc9FAd8/zGjc7/KPU6ClXNqMN
Kwbip6JCm3+PhfJdgs+n5G3rCnY15xAZ5n3wnrMCj1odr5HkZ0vBgxc3XTBxaIU5KJsg2L3vyMEi
n2EeH3dhV9/GlGphfAXCuh/IIBI6IdcbRECYapatk85UHGuB0Z3J7qM/8y8to+9UN22v65QB5DU2
00jFtd4v/ZgaXyIH2HwN6THoyxmohfEYA/6U3Wq94fmvfe5iRwegwy3AdR6pTZGqG9iWRkprLo6Y
3WQQ/GN5G9PNPgHFKOus2yyHMBYA05Z8wVFLz6Yrmypx9eR3cnGQ2RmkDG8riWOXh+FGOcvOrsNE
6KgTkxp22JxWDig5ehKUiUaZ02xb1cG71lzBIILeXNgSR5PCE2Nx2HU2UX9OcNY52fsFc5xFM8Ko
z+d8WdO4UnVnS47ImCtMOA+BtIvHItNGf6YRuK8pY9oA2T88QDSawJ55wgB3k5snBxgW4Z4Kkqr3
9CUzF0rp1MTE+WPXWOSOcoLYKFhec8M4w0ibkrdFM3nwtHILRQGkkTWSaGdGsMkVdlgJUk3yzpL9
v3JUt+dtn8WGPqr+7qqGltO5EdbB+eiTTQVsJnzFCFEcdZ/gkdoyYim/dh1D/ggqUs1KNOPSfd15
Kd8Hw5WELLbY9ZelB4Rbq0YKkhsJYQlGQ5AnpekrCUAMVbaF8Rsd1QESf6lwqn7ZDWMfsuW9i8TB
c4pHzI9oBwA+fbUdm4Hul4MCZR3zHK1g4r8kEEs9CGSblg/T7ioDKFW6Ze0dP3g3xASsWdT/tnHp
XJ1UW+v19WiTxkge3AFRVb46o84jwKq6B8vGX2rDuafpfp1dMRarMLEgoa2kxPqBI+P4MUry6U1X
sgycBJTP/9wq94XgJ4jFQVHIW/BWsu0CjSh0/oL8gF5fwk/kAzep+io9++kZm33rt7dYl7zQB1Ak
fXDWBAxOm5+gBxlksAyyv6o2Oncs/2IVzPvSB4WPoQXN3hOVniHv6TlV18UiGQD4HdA1QULqa0Oc
EzRILYqIUfdxe4sRcdGdWsfYA1oeJNbu03mQdQnlCqvjjXJTBJDNZHtW9WauYp21O1Xg1d/rJt7c
O9+56YUOOdsrywNR/zTKV/9BB+Wrur7Hqtb1UXJQvKqeS5JRvyQTs+3+PP/yvOZmoxxLIYz67ZZO
iJiEeAyIb8n/a4oCnd1yVdS4BYgzz5QDxp2CjW5L+eza3y5ERT+QyulWvUnYnJAv9I9+dd7BLzHk
ZmwoIStgcdt5giJN4bVJLqj1ItjWlWrcchgjO2szrA6ZsBHu9ipVDZ1Y+tdQFH/bfLBIH45W2+SW
8OWFn2yl9a0wm+arWHwIuL6wgZ0mjcKwf6+GlL6vHG1EUmEfpLCiYZhTt8NmrZaIN/xi805VaRJW
MWmnQNKOHDOrty2ZnflCD78NCau6PnpAusKqB0/7Tqc0dSaUkXpA5JRejObk4W5iGKXaUURb24RO
Rbpgp6K9zewsRjQujL6ZMLsXYYv7G4dz9mcuCGQHdalUGdWTDhJ64w0u6Y+Kzogsg4ph09JgNqgv
7T6+46QPZsZFricau09P6Qn9Vm2oX2RYJEMpY9VlKb8RkayA5gIV8SIUOl4fr0Dkt0djLsXVJTNe
YL5B/rBH91M9Y1VQfKrGQKge+M/TiTADnQNMRyJiIYJPoaKZtl2kDJWhzv4Tihf22FfBgP+UMTmI
hbBRdbEsP3mEw5ia1GP9rLCmxZFLa2vDaZLOvVrlIVUaPkAxU06cB4UQFbSO9tD0wkM+cAa26UUn
n9LxX1sLdB+5BvUPJ/39bxeQlmuhOK4DpZheHBZdA2nVd94tgyq7q+5AIujCqY45Gon8Un4cohj8
I7KZhxnTNON60FM7Gap4vBgyV67eA9SbyZ57w7E6D+FP8ln7xUaRrddkrfiDz+EIOeVK2wO2pdno
J15qXrPbdNKoMECLe7v3uJ4CCTU6U8IA9kgAYBPH+pZ5USPwszJiwozff5ET1CmuUz2H3i4bd7E+
pyfJ6rt7RAFEBetgbwFP3gjBpqnP1YI8+8uww2Eup/qfF1tMlrVbbPrA2+v08tFsDRxqDOMn5z3e
U998hXRvAXB4gOgjWTCcFDDlbHUPBP+CEDazLFrKL5YGppKOdsnGXjFTCPwUjKgTbWygS4mTaVEH
JI8o0M//2ndw/dlidJ53PA8XDAFOu839tkkTS+llFaYNZpdN7qsixh0lkbbhcR5hjlk+G9g4YXOv
C11bS5FIZyRs2CCwc8U7YSn3jfL++xl17Gsdf1GkBOJ7TrAa2ZST7g4a2z3wjYOkA6UN1kOzweuT
SuxuT8htjqQL9utaRKrPgJbazcdJDG8QK0N+8BYotuBWL6WQB1GBqRsoryrSxCWMZR2u2c19j0sW
q8kJnH/pZNimGGbLM+3B990aQLQ0ApQB74VHX8+kWviGEYBtwxMMJjbt3NyGATkl0zKGqf7S2mca
wEpZMaZmtI/c2Aohwr8WK21DiJwjc6XOJwIhm+gJe7yAeBlqUROjsU88sKRKyOR05SketAnJ+npc
F3JUf7nKZVwLn7GveLc6PqdqeTySDGeb8nEX72Ro3+tQI9FyHzDXZS/qxKFdR/LkZt7pEIG0adOE
HItgjsWM3EBsCaP4VH8hWMGR3tgwFQhFmu0wjv0Ba4jTSecOZ2t+4k/AlyHcObT3vVSXktnQX2co
RLeEq75sDbaNOc2kERITJqM8pnxdNHTrzEmAFYf4qPNwxbwbHnLSVitu5PVWnAezk6+qY3DlSIZ9
j4jX1l20147+TpHus/FG33oJlaGwhm0k0R5RrBBY4ZT3CHKDlYUMxVuBmAqFd1bXjYEgaX2V9gdh
fcW7JRXUKn9dSSrAqusyVGZia7iOCePeV5hevp6e0pg3GChepPUxccqEGG1BMzAOXb+pTdkS8LUX
Jwf1XG7zIS3y6XF2COWrbAS22rQyuSHX/rlbxwQjc8LUI8Ih8MvtHN+l956V9phzAOr1sX8JSEGZ
UNt5evxIB+EQBSD8GGmabEaUxvg0zTt53l2Bjtp/jHVNkRciVtgQ0IKSJ6SEydAtBdoHU1WBSzm1
YJCSd8KydBo2nGrDKnr2sQuG922Zh4c9f0Rr/JelnpRBH8dJRRcLQ35yMBMEFSZiW44rrngHagX5
KWZV14Co9hclK+KzaMF/BB0uu84HR0KEJin/x86pz5sYz7DsIXn4N4e1UqvJftx4NvLMd8ljnD1e
WFLWk6v6atsc4gQNaKy4uyYA8+L/69DpSmdNi/K7ffKPDdckI4CCSOZhBPyXRwLjT29EkJJsuglf
hhJop56FMwxyWHxzPYJPpNmKC22QmFk9+8QtJ4T7wN5dQiNhMyat8q79RszxNg/5194mZXrDrbF+
DzDL2+GA6bTWaKzxv+mk7//8ueTTUbgDU4J2zYJXzKMUDDtYIyaddVq3zMyvAYr6aCDXw+g6zxyM
Rza1T0TGE4WBpqFMVTV27CUyy+wdmVixV8VbfA4+4VnJDkzXdHtSqICi6KmVsnF8VyzKWn4Uasky
7/wr7g7jaCWmJckBNINgAvc/w+fxagY1gbNCV+nfIrIKElJXU8MER309uZGK2Ms+c+B8G4DGynv3
rxTgKJVffkzVWk/3eIZ3kfuXp+MuphCOnxZujerrVtK7CVkh9mMzua1h8454d/y3XZxIKxj2Arhz
3CPZ5RWVfxSNO5+vSp24hY+9p5GfAeMZW3xC7woTCcjqlrvhwXVbDkbYl5FROEt14c9jIkpTgOb4
vWhqY5v/h8vl4X/Nh8pR4QxZu2G3JwqH150/SB14L9yww06ZG+k5mBEA7Ks6TfJzquLpE0/hKxvG
KT8ay4mCax9ek5qI6Xhp5W39Pr0r1TYCbxiTXNrBGtK9ihf1hpBJpbd5Zj9qZVvXzY93qISbQqSe
Yk/wnhQ1r2QetgB+G09+H3COCrB0y+ikE6gy/+469L7pNHVraWcCWde5RQc6BQlJTT8J7hJnd82N
togN5L6KzQSiVip796ly4SvKKzN0SY+DGeRdKQx8StT5y1kqlo/UxqgzxYN1yF1wqeVi8q+l5usv
kiI8JnnwM2gRFE/PM4cq+wAMEcNz6WWdCDoSMCSdnUqIWf6TG8AV6grYwMCm2bOvOesA2KuLMmwv
kseGrVHBDYMNsq4bqgXSsra7jA4foXU/UDr99kKO8UNRakO6Or/EZj41aIlLN9fseYpjL1WawclI
iginuYS3tM6SDXHeos1w5tZmonjW5Mo8uK9glA7u2M7Ad+mBt0NvRLf4M4j9a4WJrjdMCXIYOyFx
OGbqM6R6kw3Z4rxy198v9OaCwkwafrPRvp2pWzkkKrPI4QAtVKMBeeA8UBoE7MSbTRasTOleGZ0U
6RmEtvRTXSty0FYpwbIc/Mf5DWUMAoVRlWXM2uqahph4X8nBvNFz8dkaHTSjYTRypjFMUV+m2WBI
wA4AItp4ABXHUjQ4T29KXN7KSG2FZrcQ9Dmt1pvxnW/cfM9atijORZZL1tQ2cccxhnqTns3KAFxz
q6f6hg82rS9gUFCRGEEO8he+WIddSV+ZofwoYLg9PUHiYi085p4AvunrzSuyx9v33Ie/pqKe3grp
Sq0qHDNjCVfsbkT0YiT44N9e/uzE/cQB3u/R6f1Ydl0kANxaDaqkTC6ImnLdsDGVOUH7qk0/1ukw
TpdIJ+ArK+I0Todi5BnnuRYXpsXiCfdDliZR2KdJ2s/qJ+tnlh9HzfWLHzk7p7zx9lu1RS4ZRluz
p/Fw/3xML6mZdIXE3pQNZyoQN2rsrwq63+wQ7sJZlNBXObRkIhgwVAfaQfZtYv6hzNT7g3+mG6rC
SGR47J4tFteDNik1aPxSrNGeKhfYjGZ7ID44xLkpSQoIntxouKnJgQw/wtvKXu5WG/9pErfiIg7n
NAN1cWPepgKs1C97bLqzuzpSOfwZwSKKrcmq6kh6pH1nOuN0qcNPltg9pAGRo+MQPaiPyManku3l
v+/i9R6MuoefVkvkSyNPM1+MkWgihmhxOGDBxHYZ2cxl9XNYiOzd+U3d29rRSFhxx9C8M7O1Jn+A
4rlT+A7x4UoMDJd/L0sFGeaCl0Fn507X3ePfwTgT6LAA/85qF7rbo2BDCiEIRJUAwk/6BnL6vYOd
BmQNRVOx9OB0amEjd2Kp3fgmnBWG9H2a03mpOm7cFiPPiDvlYcsiZ7t+ifaQG1MBUf3Viw3PIaCV
ycj2vkHULX6hqoJRrsRmW/jcBdAuDl82l7GiOOAgEBfqdc717efzqudQ/SEnw3vHAqUJ7vvF413a
l52Z+8IWbTTsZRZ94a1oMvhQDsFs8be72p8QCPSKj7HfBmgWYwvQFYFogUrbdoJPyKy4G99BEJrv
9lZX5Vu1InG8etN+EfYo2fNr3KtO+RlHzSO+bOK5xyqFyn9+U/va3dRLGp67mhLT2Sa3k5LyRnYm
AhIajnbQD+ZBKA3iDTgrCEdxRyHPB0SQ65AyqXV3g+yZJqjJB+WR3X3Jl+yWK64wMLMfoBHC8acd
s+DESH5Z9d97zIVfdqJobKFkw3cXsftq3rvV3RdBo9tC684iAShq6qX1bEPCtdCJI+/yVnof1naI
vUQ7uji3DMqNx0l7+5j7ttL7LikHCob71sOFOjISZl/ynHWrN4ZRXHi8lywF3GNgNwmZ/rCslewn
5U1VC1GwRcIBmlR78Gw3mFbHZLbomWr7ujksr/+PodMcKnX24CphZQ4zcUatnPZXnlMQQRpRhXxL
PxL4NUcTRg0jGMnDJhF9sHuzwoDPk7QtqinF9iF+IsYTjGmGNA4Msd4T1bvkvzukVJPI0LLR8xuz
OIgwnt53IBt/iv9M3jAHZ2Z5vyeP5jrsRXYU8myfIZuGB6y8+9GMZtox+6Zi+VxESeQwHlfbIrAm
Vo+xv9RKkN5QWOt6GLElC2iUsYVrbhfA8bcX/7HVq6KXJedbBXS76uI2Kme//OpdFYq1pdxL4msS
/xcpELvXbTMjyDetuEu9sVOmnEa0Hk8dagjUGTT4eBYjpAqr2W13x6GrP2ounVFmcik/8y7f18k2
c9C7iXos2ei994cDfcDEh3rDssDlwKDuxRr0uGcnZSySJVKRK+C9sMsGaRfTnXUOGQRJo1lwA2p9
SwJpBhTEzEu4sG2TLMt/0XgCfbX8EY8GKg2zyUdLX8KM3sQXc2BoK/BiWmoVlU+WtwxQYEy2iBWG
8/DqcjksRag4cqSEXQYJ5Zdp37IJFgqDAOBGbTbGcSf3/1bU5PcmLFx1hsEHpX9pXvdfcCa3ti08
9gs7lZdkykEszolTjKOfiUmS8XU9BcCmOPZ2mAqXdDBm4oHvimWcOue7Q1+HgpLJxnYGdhoNRwQm
iVrmHVbJkCuqY81vgkb6RJZHnL6XdLejibXfGZLmVCif2yTlBfvB7WgRVvqeBIPpShblBV0fQmIR
REi2/QpgFVaxcvI2+vHvYB08XfDLoAY/nO2LrgIRQ5ft2fkywDrP3z+4fdgDF1sLojxLODjSRMzG
F0r29D0Hl8UTIjaXTyvqYYyAZE9MFiQoMi+DBgdo8LWgHZeH4aZwi5f4SWWMx7dbVoGL1yu6r7N0
JU1D3ztD5n/Jdc4qZuFbNoQWg9J1Mk9lGcgPWliQJSKWm48KI+9t9Eh8ToZesm5QRbZ9SPJxyaQM
J6GE2xCfMJMCIcemdzRvVmHNbu1A2eJLkZgWwnRVwh+qguSOgkgnGD+fz61iSxkjXqoD3FK/7mxk
Vru4MIceyG4VXFtuETnUGqLgbmyh1TfLq3lXwnSJ286GMBGIYFA3Emy6eeWbFMAvRO0cFlwirFW8
f6m6ouLUZAC6ktDzNpcOden9ZoslEgnNSkoKVCUiyOiFueFrKAnOmlB40LeTYnVxSM5szB8w+R/R
ST3a+0VWuSZ3hzR0oAERKGy+4X+gt282N2im/D7w/ZWROe6+U8wG35t6nFNAZ8Md5YHqqP+uflMy
NLDFHhHwBHyIEm6yZWZSVrN+2kXBk986gkEPL/kSINDZr0rRuNSUcXKx0F8tfhUh7hk5rdifRhXG
atyE8kjTBXxbtZo1igQmyBfYXcF3VZgBRBwt/nVf9+cLiNCn59IMnb3exxi3MMkDg6Oy4IndGQ34
jXR+hK+KWKEHCrJ0pZZgPa7aY6eF9Ydbv2HVdvAw5wisWoDs/5BslY1CWLqxPXuds1MwJohQsZI9
Cr7C4gq5utMjQ49Ct/Ovldw+8CYVUkwVpIu1bw540d4MqinpS1bH8HhcdXgpMpWvMC4ZIQdJiB6n
YJ+GZqPt6sbMsMgVvMvjIlGLW2z6ENe0plJa5/1zPY4IV9weFCds0nJecoM+3Fcc/xS7Fub2Sf20
ixMnYYZbsokViS6FG6DjbjKrNOd5Lbo/TVMaLt0aOR4/E4L37vBK/S5jgBIN32BQfwBNyBE9gTOr
L2AnC0IUSSg6z3+ogeJAuk0i15l7716zNiytChyJI9u0I0TLZizedplnVvuAX0iCOisyrqCkzZy/
JXWdVkVvxZrBQJ8uTBmfgQGou3zOo3w0HnmXDs45eAezWK0NvYOpiBOtH3hg+nsajTKZEyoz1QMG
32ZFyOAgAqY6zEbQkNhy0OUPfrJKYIzDzl0uIlcG16dD2E3dvTO8Lp9MKAtokPhya+bbLeWcRmZp
/4lNtsciS3gvYm/Pc6paopqzm6iUj+xtvWTgBFEUyHvGiU9r0SNyYxRdEQPetcr5l5TD+ZfI87Gn
IwiPzdO7Y4fnn/bmZOJsgSy1SREgDymi53Ywt9jpBsJqHe0RY3G2QjU6V4E9OxUvsEHkqARP+Wyn
JUTA7dGSjoLGRPFMuNig15Sh9SrHY9/FfggjvXhcFPJEwFKaBXHuBKAueymDiMcRFctasl7oiuzn
l4BzPvXE1WbCxuA89VGxTFxhC/de3TtwMNYuWMGDLke8SbRA7j+88ugjzeu7EIbv4SOL16zlTwj4
u4mVkOXcFNxoIVAp794r29QTpIg+9tnredBACmbaZjTxRqCt2yqGdjM58Ic9as+vwFONlbM6s+LH
kygVOGWq+LShywgzGGjbZNLO8hYKpU+avAbufPTPR7CBG361GUbqK15fX4Px5x/JmRb4PHGeCggX
nzuWfTVQpQszv+HpuDcvQNqoZQjA6E+QkwdI2FfrFwAAyfDKb0/gSEqNCydzBIL+RzzlH+JFuQv9
HZOSIPl6xrruZ5E3cW8o1tnPu2tG4v22hRzoyEFcr0/GctEgLQB7zLSZLZxAdFo5Jh2a/9Q2Zpxd
pwu0yxhco5ZhMIPVkboL85qvQuKl9y6TgXF5AJIkmVJ4BUrRDlnQcIaGUAUGqeIws7Gomvzi65gD
yncezPwShXTLW7dDhaYU7b4qbC3ihVheRdtKTPmaB+1dgqc3AiSkz5ge4T6qHcd6WGcRTLsoZrrD
7f3iVNjVhXr2zUc6nnCe1EgyE/1wnYHEWFvUNUO2dZOganEH9Ce+PEpRjicJLOL+9ObuOZPUB88L
b3L1FCH+gretyzcpj78G9mylGUAB9MH87OLTmmgNZYMxaXxxcN1RTemN2x7l+ilgRhLGlD2sK1SC
zXDQ4qGojZUWzFEPU9SGjf5Pke7aUMy0FpbWzYwmGA6zCkKITfMmAznYxBe128PogiruQaibHcO7
saz0DZ9y+++kI/isO0RxUrtTBTUV2fDRWnS/sfAaRqTa5BlkI43XZUkPHw9MJF3LR9F04HkNJBUf
ArbBRRRImxvGIUB6X0dNuLJxuxakpmrLwc/XKXb7f2J92ZLw+/WKLDJiqm8XUPoHC1J1y3LH4tiU
0XhDPGjFVdA5h1QPBBNbgaq5LeX5LiZox/E8Xh2Vd+ZmJFqtrjWTtQTirayHJQl55QWsEWuHrw6/
o/BJhP9arxls7REfN97EwVyWtWFfQWXLSURtM7Rzrba9x0DbyJOCjz6sLqePk32BYxq3ZliqzvcT
LjSS3vDwfLHgijeuc4hHGsB2iDWFrjliR27pwcwkwdok91QpHcNJe7+pG/jSUUjBpfWQJWQ2OTZg
/38hzFBeww2yT0znEnoheQ0PtqnhbphTkzk4wPOeVRWzk2YlEkMYt/NwT87Cfg45OAZWyZ+mAYeu
+V8WX29qhee3g+J1g9ao/VT4uujGLFlOzmiRydFf90oS1AE2Z91Qc8dbXtQ4qrQjOy5cdyXjoJsa
92GSTrzbc9xjD7olauR0YduuGot4IIZU0WzMlxP+YFj5mwAl4N6YuZ9x0loNuAtRLlUrF909ur+l
TJVWU/EadLW7jMYOnQufOZbnMnm8um0tANKwtuj0Fmb9UR3IeSlUcsjKziez5vexJVswYGRhzOkN
p81iTC577Iqvj0Cs17RUJdjeNzw3rygOJ6ou9B+zot0fTm8gh/XviLuSb6J5rAky4nHMdmi/uOx5
HWpFU4Ad5bWk4M2WIwOD34nVOpXMI1iKKogWC491kVi/DWGk1uNj5IMiWyRXQ+iVn2UMQoFN674w
D7ysK4hvt4/SDEmWd0ecWC2Od/HCAbdc5M7fNFakCAnsYfjJH3BK9DG5//du2hwTdKqfZUcBEata
BuI9OaxuNyOyrxwicJJMtNgv2m/haRAuQOeais3Oxd/0ME6yn7Md7YpYQZ24OVgGE42YPzY2G3+A
fDZIV/jQ8QJVgGxNU3PPNXFflOirVne3TxvvdwzIQDEYVfHFE0Fd9EaYs0nS8XhfLVUKLn1HiwXW
bLwlv7QmeVL8EbADbP/zCYp4z5E0vjD1VX8AMOLP1OWvKjykq6YaG5VjK2nyHBwL1n/jQhQ6MhIO
nHkCXCR3YZRlXDUpNFDQYPRkuevuoG9Vw3tfp5/i7/F7iL4YhCAmsxnRb/IU6rTZimMPb8PDGITL
4IMBP0kfADgmVs65RgpIfok+T7zr+EPN+nV5eVGf7e7o26ILKVP/Wu/WdU44cu/XKKu8xqZw6zS0
55UQvcUZRtnRAJf3pLQIaP7XbvnQPzchu/9FRkjr6tv2/KbhIz25PlnGY5WTaEDGRbk+IG9Yls5G
95KIddEPCDzBdaGQpIvUW/LWOaaQtGbyo8GaFMQcp0cmjgs1xGOiv+wTy8qXiGZgGBHrBHhYct40
aOgpDbo2H4fDYRpQ5WjXeYguEKUi6Ab/MlBCKk+lvCAzcX2kVQsDQkUbTq2xQgDq74tpXujLcYzp
t0tJSzfwYP1k/vLky3jQ9fYG2ucwke4tCabgqA/AUObgtFDMJmVCPTcJkPc16s5FiCcyv8ZTSvZP
9gFMXH7lLyyx2lS4bvtjnfPr84Qi9Az1Dqc/L3/qWBLEEwGmo0e4Hyy3T7k+3Ufg6AGkOVEOXsgW
3yxUUwhNVkRxidT5v/ckxUbWdjwOnE+mOTvLPtRIEo5GsFUr5rN33A9/SCFNAecxLySsZw6avEOp
vwCLUqLOa6tP4p94U00vTXTw2kuMuuZSHNk25iRMvtrCDwOMxNFuZdD2GZJeZx32hSY332TWG12K
zXCuQgOcKP1BP9xfJ9dru27rS3wjvz/MXBwJJCcXWAIwDu/GY+Xm69L0/1n40lpR1a1A3mPJaFMV
8Dvw4Bqd8+00u3yIfzlzbPuBpf75hwkzEXnhhQOPLtm1gRPmzEQIizPZvjEhrpZTEOTVNPdQ3w6Q
iSyttB/iBYawxqenVODH5rBpVL/a5Y0Uy9io51YGZl/M/FwDA+SLgLutolNRRgkHXtahEXL2HTTP
e+9vxUccyk/om+xeRGPW5imnxdUY5q1WSjSv48XqjOP65EWo0KtK0NAgeQ1y9pSnoWtgSss+Hywj
MQj8qqPN7z6SpBHNvRkEmCAJKcixx6isDaX1Kd9uRbbjXDwXBQiIlcm+kKLdlkpIvxeM+d9iqeUi
7KowJ3s0S4rnfAqjaLgCZy3q5wyx0h5l4KpXaHcYsULvpxdgNrDypnX0Dz4I575X6fH7PEFKTf4t
cQs3fgTbdw7u4gYej/Ha5yd9MysnND9yVW7vjqmxFCOEbnqHxrwU5A+wp07uAIe0l9PTnXrS796D
MR4/fXLIpGJ1OZlDuaqEgKDuXDlk/8u9Im6B5dC9kTvUz9Fu/QsRnur14kim5oRpRzi/+v0Dsro+
LuA7WKXFnXXO9HhhIcMlAXV6W5C/lVFMiwmvHPB3c6+/yQpLbNDMLQs0ufOKz6OJyzUC6MXoBFIY
YOuJPSh4A7bBeWf7LuVzAMagTL0BZV6Cz9y7oyB+Jp5sqROrZEdoZhIDoC9PHkEFlHf5hod4nzM0
Y23ILEl+yciQts+LUbRmRjOUkE0mQRgg5rXOG5gUSNrJEr1hKTz9T2J3M0EGpnsYuBJCz0yPLgSi
5qvLRx5GZduz+s76o3f/IuWsuGvc2CCtQsIScudOANVdyxWtxyysan/759HImFGY9RSsI7behmSe
TCEaxSWFjo25FbF/PMo6uqr/X72U9wmWv338cWoZSXkTAcmGtTMoNDhqDwqK4ZBDyDiBwFIjzAab
cMiQ1S/sGGv1FqnyxMRHzxcq9YGgnEcyy0e40A5wnwFVpCKPpqyVwHqPOjwLuz3qViyJ8Nv39gjI
eoL1Fo4pUDXHu6I3DUJQWIIN12PAuyXXn+pazXqRMk9CrFeqhULYP3KO6nsCdj1DYideMw5/lkLD
9wAJAnZj5sSmoZemrn3y+vk4Athp137WiXNGNqSjm/sIeNnLJqi4FnI52ezxv0PKFjGsEiN+nkSK
wH1Ivm5DclYdFwOu5A7Cva06gR4qtbEgyN7dwhSie7UP6fFcqaLZp58QcpjFW4YhgtSAibpvDax5
bN+xK55b5/E1vcB43mHaSfI+5aZ4RcK1gD/EXQggpVPS/wYOynkfcLAXv78NXM+H+rkWWqcaZxNn
Dam6qQWUIGnGRmWLnPy20mcNWyoewjBmS0LdreZtpm6cr/PHn5e+2JkGp0u0JZRFZ3dIcIGIdLAW
bDGP/xAkpMR2u5BREtsHrjDxKVcOsWIdfOCttS8xss6IgIY9wRiy0t7auNW0Oh9IDB6mYC51NGue
B4acm4oLNyHmPifMGRseCEdJBne6svECBEhYakmVjkbWxBG6EtPQzZHOgI9lfNtcje8wdRuk2R1e
fC8aRjxPjWZUOD+tNIWVUwhRztm8SAqmMEP3xp0qRF+7WaDjyX9nShhgbkfDcFfdoV0Aun6+PVd5
bSLEoWCkeLXF4iyEtkDPmwskTZ2l9k98LtfKlEsOIbI56MPiO5xV3jQVhzMr93hjdNQN0P4OqQnt
NGyS+tN+xZOxnQkAFx7SyysDfzGfvScByzB2YuWLOLloUsczBvD0cDtq4j2IRNj06EAMguHjhqvE
Irc5ExhXq4z3ep+oQdafKbEUXQGtWhJGcxz+eG/+0E3ZZnIpoJZ/8QumQwzKBdbq0LE//ztENsvQ
N6t1eZE5YzCHN0J/QtHcGvQUSD+bssDHosfoJ14yqDGprrRPMrPXw/70FQpBrtG6bZxcJkQCsvET
ho8eyBiYzUGQz5okG8SElSNIrn9vlCIWp/DoiCeOdHJKHPTvaGhdtxMe1PV9VSB916R6WYI2+2rY
XR+koEoRtEjS7Kxe7kJJ4lBw2vpab0hD8GfRspCtMsVxECcBDSknuTrb1/+quDWOz2MR0kJxL0yr
mfIkXRVfRMzKlGt3q2Ml/We3z4y/IlY49uSj+R47NL30+IJQolJFimOQtoP6x7wLRer1jKGkR34q
AsvM4bVB7pMrZgKMUDdlLMe0TdV4zTo+e51SgiGctlw9zdPxRUu7ESojeoTDG+TEmcY0qISbFDjr
Rcwzk4aAu1zrFYCi99p7PxUys98+80+KXupb2TQitm3WTo5FzgKMSRkwwCXUvXUTDcUBMDKGS3p+
f1vcOEfHPSdEc4noCrWPErsr2PhXlzrRjRD4OC4iSPWqD/q1dHq5/2owsD1LPgv1QLHdPExTz0oY
pkolcnaUR76SfiDFM85eJnx7hIBzU8HJLtDVZBAbiaxpq1JpqUtIrzW34kFFK/7qPMS5r+rpZaXD
MqkCmC/2az2qr6bmuOKiEZbXDU9Vtw0jsXcRocJgj9YBhIzfmOfpU1OWM0jHrqa8NAK2vDprBJ9q
lQKM64kaupzgkgPGencGyf2FjaMBU1hBYE2ft5DG//+t9YO5NwoCCYwdjM3cjBZ22/yislBPTpbX
b4qcm+I14a9piUqCP1Aat0OVET46ZurpnGyS+7hjfCfknc80UTDmPOPGSI6tqWctIuMzgympwZmQ
TbwGjGUI+NWdzwwLUYIuZkBUdfd6Uwr/rtQt3QRff6NWwtrZq+fuoeJ5C/kx0J4kC8C2aahHSwX7
j+dxK4PdPJwzB34/6ttWOQsmLi2dTjkZJF1ewi+4F74UYqbBnnsMHXgdtk4wUIwRj5W8F6Yt8lx3
2f1WbXyB+frMaYocjfK4qWkSp+gdzf2sZoC2OTMGNt4Dya9BfKLKWmg81PruqJQqmhvNjEitUcvB
1YUtS35d/cQkj4e4ySqppuEgvL5NFhjSZMMSQXHM+ZqF7pjq7FVRiOgKXDNsXgvvWZIgGvKrCX50
iOm8xBnkVfebUto3VU9WuCMQg9MgmmyrPqKsDSbQxAW+vKiJBvBQ6kuKowL9+/6nPasw+mf4L4ug
nyuMeJs7umIQ6TzYnDbZ8rtYfqrqCCU/lZrokg64A9zTWpnJ7mu+tOH8PO+kR7YvMqsnyPVOkqYL
VRcBvu2wCsJnoUNXe9UVlh5j/+cLCbQlOhn5TkqRgluxxntGGV7A2bbRGrcyyOdBg36h6YSzgnJr
dkaTBJCvtVg9C00XWs85FBaIbADMLQi3EZTfDuiNeCic3nFS43NUO6X67HuKrnLy5fXHcBiOURpi
Y8MCGOxeZiZGPBySycSvscnxk2YpeWeXXmSgVCZRBVni2A/+PzjuudJBMCZIfLbG+Ov+P8G7BGVs
QIwW1Ixa+I38y/JNfFQDeem5ddItC40L/XKq/DL5NSmSiRNR6PAf4eOyquOMwg7mPoJAil/G8FOO
03o7Yn4qrb58+gVlQq4zAhFg9es+35CmUuQi+x/dFK35wvkctJYUV4LN5NuLwRuhjO0+rLQd9HvN
7gGhkLywvA5iIhTPtuQyvmZ1hJPp8/OGDk1pWzq6nshyKLpvD8dTlJ6ZbNGnOBNG+KC5vXQgLCG7
M687n/4Stdc2Rw2S7PR9OpVdFBs/G7Zk4eCIv7rF3yx2sTPzZU0qSmcskw4oWocY5xOFMP01hQCn
P/BkmjtENZT1vKkp8TWf+ebHyI2gyDUx7xHhgTvCfNGycx7JUFd/NCqQeiooVGMXm7U4wNfcuecJ
/+mFApzcXZc712IPOMfKxiTt1hWmB1DkJj/jftlXbVUGJe+8cIEWaEIOc5icFCJ2q70mo24G5Hh+
zMqiZGp8ncI7AdZdB57aeNC0SowA/oo8bHPNMkbWh7yZrsva3byZSpW2GYsXhYHNC/4y3drkiwrJ
z/wBmxJXK6e/YcYYEhV8bAI0YcF6BvPDoYg83dDQPLdV2yBzZfdcrrKQXUq01sGe2nS3P9yuFP0w
ob5loZ8SCHXx8jq37XPPtXWxtF7rdI5tq0dfdGBv7wvg3h57YF8E7p4RqAI/IeaDnjscggDXrjoF
Mg4Dk4vpVVU8QyqJI/nyf7LMyLdSZxptrAo55e9yesOJfhZaVCo4kZTBVraN7rKiNRgEbWd1t7R0
jUwg0GdEw2nu4icbUUrXX3ExDmdEyQ3uephXTDRB68kzsCQD3gkuO0gxXZCqJyR+kX2oK+Gjs/me
tHI4lkHOAKdjKWVctM61AkULb48Zc8i/hMSPJSf4qu3zXbWvyxpCzehJUUIL4YnKYAnxzU/3PcEy
NfcEmXknOmTX8daM/PWHMvyTZPY/uGf4nPuhd2F2MVXVraor/iKCa4CT33tUQYgKZZmjYrBjtd+i
3uu85N8wcWsRxV24ZANTHCNE/CPkUMGDIMQhN3tB0Vf6V+Bn37XEqqQk6PS75Rt91uM2hRSmGmHW
70mvg8+UkEOtejKe3OSvIRUqqPfpRGH6xnel+vY79EkgCjd86Cz0+g4az9zH9x1uzsFq6/UGKVek
KYw3x83qIh1zYBU/+/G0h/AFdB4DhUFnbCLV0U5zrfdNFp8nndQnki0N9w7oLSk8mw5GDP7udr6O
4UHLaFE3KZ7itvJU/H8shzwEJUcPNCBYBuwsDIXsIrVjH/wOMtAmvLzhH9pnIcbAN8+kJ6FbZyjy
FCNWiEDrWfodN4cMdDZF8FBld+UlvGs3fygq0/B5sEd3xzBB/uUtZdqPMWZ11j6YXPqk+fF2whP6
vOs8vp6sXQOVknRaLZTKW5Y8oDX5m0CgTqovqltUtiai9na2rO1dnEon9Y+nXIIfo+zKGdzDcZjX
9Mb6N2n68i2dBrqk36GM5qVIhgcC1qzth6J1fRDn1Qa2WSBA8u4LNiqFyD0aSQErIQwJdFTl6bje
Ng7I6GIAQSCntOfJGE9HQnFxg3l9mDB1enRfcUhcQGWfOVzhnO2z7Rks0/nXTKCfkW/7AUKHEMRJ
I0oSf8shS7eP2GUEl+yFx5oCHigJALUT9qd5Qj69WtaRN3fjVkObJxnZkaMwhjem+hDjNjrUKQtZ
3acpvySdRYYoq+eIUKojw7GNOyC6el8zFPLcqdgRopXnwHttJyFOMaxySqS8qqRjHzDi66WyG/Zq
i3Uu8CWU5zDDDSJLNruArKUHzv3KPMyZ1Ktttcuyq2/a12Bxb6d7HK02Z1LSgCwCuT6vPgYRgS8A
kzEI9yV2Sl6syHMVKJLJHiv9OMyax+ttNgtw5vm+ssSNrPhGsugvULwx7EFUHBkd0UDvFNHtLrev
GMfvtl9v1QFCJIUSi3O3R5bsVKFCsSnXcHQbahzDDkk+Tulc+WPvH71srRkaDM+JE9D816TJ1zmT
504MC9NK9qWgFpyOJILVfW6g7o0rC+NKVgPsvTqQ9LJTLNRmsJV+g7OjW1yqdN8Fw+Vb1x6gT+mg
sijnGwqkxNlVLNWjc843e0rRfAxIIQER+ngOQFW9Wrj0LhnBjAhd/wsrzV47fmgd50zjHjeswVsX
BZN9sZjdVssMwTnVoYLWi0ygYLVgsKkGZyNFY5FenIJzTImVZQUs1uJFTBzWrQu5yIq0iR+atkxb
tPpH9uIA+XXZeqkas/5a2RBnyBiiJHg3+LSJUPYI5jABKQanICcXsSTmEnlUxIumnvZxdiYi5IwW
LELsBx2TTf8Vt8NjJ4Pmej1RpM5UGyVq0g1zRkTPW9X+u9DND7gNchnj4DNRl5BtXA1OG+29112t
M3A9hcB1UTKMUpOjrP/TZC4qBH1qAH54ZMqpk4ifHoVabGlwSiCpzgJqlkj106DgUp7IG9zAaFHh
LQCS1g4NCw4yMYtY+LM4h1jOb0mqGEHDYrmdIcl8zoRWr5qnWrNX6oZhk5IsKSuKYmGmcBStyclg
cRCqTlzDU65z8yqi9wq4L9EWUrfHifzdsaJsojjefjqDR2VTAdrtLiDyaJdzJzbAFLPkddwpCVcv
qijbz0UqBgUOJ3/kWun4xAU9oOpqNYY5o41uA3pi2X5UQSSH3pGnl8ys27/kzL7U3BpG/8dTZ02v
xlav4ys3/1jnS9k0MYEksxKuCbXYrdGAucc2BM8QOZx2vi7Wzp0LMiKWXUYeNJi1APd7SHs6cKjd
4tmoBOqxKYZ5YlohlQt/e4AqiriDLwDkYAo4f8ZLhytOxprhqytMsx/00ZMxY9rhDIlUmN6UW/7y
EQZvlDOGyk33hOg9Z4uApSiQ7IOyhGfRQBa4JCIj2sBXOYuC8bX2YCMtEWoLjvbXcQCIkRN3JGRX
goG8MrSI4N1L/v/sgY4bf7IXymzYeTlg9qzkSIH7HhfVJvPx+9MOrNMNEuqB8YeBJEjVHGYIeg9b
dYuuEnYwbGTqXxI94Ym3LAwruJkx8peh5bJKr4gJ9einZkUN7UBZSa5tA4MDX5zE/Tim8cWDoH3z
PI2KORAN2DgV9ABMPeneMUH9oKsUg+OpZYfijzlLepxzTmaV/3JcyDUOKLG4T5f1HjgFTByrdn5v
Zkv2etauYrh/cjr+UUS+fTFoxAXhx35stMKQM+2WXLd+Yg4C6L061WghOnsJ5DDFBxiaCV5lymbZ
XQHBTKxFSlQTVsdhKEMrR4S2j4UKlblDEWv0J7o7IayIfJH3QjPzmNDLSF4O1kduJ78oBa/Qjzqz
JC3qNComp81kFGbZOCi1v7AZmbtF7IssQdCnM9Z/xIfUBb7Ht+IdA9X8PGa+0hMYQRJTwj799vmF
4cEtSV8s7HvXWro1z8CgCzC447smink4hdhpKCIEHhtw2CS+Ecfk0qAYPwo7npub7Lz34IFTUa52
a+5A/OnOWSAErKxMsG6/ByvnsQ86c1mimyKHmyIcRbaMjY4Vgb9JsijEaspqxy9lHT9kfTEqOgTv
utVCpbLt9ggecTBo8L2twXGRZ7eU9GVhyzDFw0jjmzuxdpqxQlRlRzHn8d8wvySNqtxVDSstHsGx
oq1vA0RPCw5MPV+a0AgQOkkG4FzeezCEh/O1GEAnmAo6Um6Zbg11G+m/X2wYsX+RL5mAtPpb33bC
SYNljWHki3guVxPPo7G5Yd46A/PC+F7+UdgeapN8F02BEWzR9ex3qks/DoUeuGQthk6y12bKRCUS
GGjcVXxir3fdEU6bIwEQjxMtjboF+JniVMyZ0mq/ZIsnWUE8fA1lDp/pwVnhRAPKUa7DlrHtIy0Q
7ABrmbQ9ZCbrMpQZ6AeTiMEIpgUcWZrjP6vSgbp2T+s/sZCCNq21cGT6znJhDldZsITFCi4FtcXr
G1FpkMEWvlw435IMthuYQ8lH35Z/ZZjAU6HjJK2sZgp//VrQsHi581uple/u9oP9vPfviLfTlG40
oBBGF5zyNmp9p0tQg+uGCuQX70He5/BJLyTjdYNZB9hioszzB0dUi64B0vCIGsodlsaNLQSE3nK6
5DgGA25KOxl3dQN/1HRAd6zKeJmg0E2KKnRYD/bCqzS74ABL9LJWTBJ4gFy4t4A+aH0ueCQNItJo
E7Nhk2vvPIiBlgHKDAu/TnW/HlHvkFMjx9sQrXTE7yHbSroT2S2buDQOq8X51ofmODaNz6pDUFdw
NUDXlIijJZnL2Za9dQfSp8htdBkeT+9FWCjN2JnKmXLx5w1V6KCC1SR4g8EzNLFNsUZF9wyK/4+W
OnnGC9FN3fKO42iWQQ+57Y7XOlHII0F7lXO9OUrAwJTVc/HggdKG1MmOVbmrwg9iVz3E8k5N7oIQ
S1lInfPnLd+A6F9aLGFBx0WCkKSK/8qBaSYOCk+yrfUB3MwtCWlN0ck+Rs24SW3jqDv5loKJrM2w
K+EA+B2HJYq21OTrZorhXTHY+TovFr7tmjV2BzkB8tGi2+Ho3Xizqaltt48Yt/eQfMntTg6I3FyT
5EHIVy8Y5zl9/jfSN3HKl0/XOymcpAeWqocd8Kz1dXmub6ax6cIV1PQFHZVBy5toN8uqrvWgbRKs
lAN63o9sUcRHueBNTGF/Drz4lGBUJAGIH7r1xR2zgFndFMsrRH7wKQZrHfCubpCG/bm73wjjY2la
14m7ksDxL1agZxkkW2of9lGMS09qYxS7IcL3+J81Zsuj7ayYWu/YhWdTrM+/gffsUMD3e9INcO4b
TkT/gVg9WgA1cbQB81UBjCwIG32U7xz/OyaZ2MHqMHHHHtjAONvAjKur4+vhsIjtW4tQjVzcSLhT
242LGkXY7HFmWk0GEkgBpMRyOReT3H7mcdvGLsU8Pfrz5SzRamQNZSxjPrV8vYnvYwSyq+kWkNg1
pQYdqszsGY3/KxQk/v3m/3mkJIFSmpG0LB19r7+0dZtDGu23LGV/HTKeaScLY7lBzJm2qX4KX8zU
/6sREp4u0ymg/jV07Ki+YW8SC7ih/q+DgAFWLAE8s29sZdSUHxG1GrzhOxGXKBmqARIr2ZGxRt1W
fuOX/tsNsd/KFzQrEXAAqLPN31UjaQc/Qa2uosG0ZOXkaTwHAl454w16rpo9Cf1c/X7RsqHyMz56
McK4DPxG7kk1PJuWZyvuwDB5IRfhv5dvjiDji63tBj7YqLTzs03BwASBs4g0JkTD+SvzcfmmK8zo
f7jVatNMs8K8eJdWeQ3iJdImkoy+w9Sqp5nqFR43yWNDBdoNP1HDtDHCPFKbPT2FWIVxj08XeBd2
IRrIQ1LpOjs13JwCVqw/14QNTu3AnGEBwv6RZY7UVa3Eli/R/c6d629hsFKLepj2heG3IbcpDrrx
yQlMGx1T429cs5FMKMi9nsYg0DOhLNduTeGcSew0LHjE94PnPUUYWmQNMs3zJjMC1+BIBiqBrRqC
As70NkneloOUL8NVxKSr2al5aGpVNnEP9m52CdjzJi0YShbvfxg3BbX7y5g0aKqNw32mgVQvGeNC
HOPX/yDsV3u5w3MyxXOhGmfJZpeOCkd9w4u3FHAejNhmj4KrAK35zI9iwJU9bylaRJdG7iIbBVWg
j3Y+W/KOMKpTOP2npV9XtjhqHh71lNx/5/jm9z90CRu5ntPDiWN0dTHDus4iiIKXwfY9zHgspIMc
wM/GoXQPt6Sr7UTLjXcwo/FiS3PyJatOYFHaE2LpODSLD5DsD6QzIThGpplf6XmDqu+4fkammcug
sLHP7qzIvZE7DhX3ul2dQHi9VhYgfZ0tnfroj164ohuEXtzsWYEiulRYCnX/jX8fr4dqevOOBDf6
ltvs0KvWXk7GbOqNzi3/qOqzUXr8MoyTea6GSuq7xa8tGpjwWPAYubglqwu1+f2nhFcZUW4qE/sm
P4D8V0R+fhb3yGzKhOgB0tE1F3lmGzO2K5WXIh9bHJvJ4TsbkCLaZ+TSVRrwTtDMD4gANPUpCR5A
Zkyh3cvCl8xJcfz5tm4q5lKd5I1oh8RaP8eV4yfWCUaL//5kyh+pk9E41PZtO4YFt/V+GPKcdAec
Sgud1cYk9jqoqb9hO+Km+T1ZFEvk+wF1ttaMAnZz4BaylWbeYcrzOjT6a6Wu3xLnWY6qtEJLjx3v
5ccCOL/qQXMpYodmQw0ZLHN9WDMBeDFGaoigYV+2CZ+a2pX2afsRxymNOShhQwrHv+/eiHUCt6PL
RYzlQTJodSFr9H/vxZYsRxJqarOG4zUxXtJfGAxcFi35cayLMlLpw8oD6cq26lIEYTuwiGL8HuJy
f7MF65xe22V+40RH+dhM6O+XZVlZrQ5GaFLixeHrJsquQ1KCdSdI/4nib8dNmAVUfy3HGQGgPpCZ
L3UvF/4S2bOzdN+1QwVQEGQ+E2mlJnoaP+vcfX+/08RnzxOBc/3YcMo1antn1Vi7/5k54StGXF/0
h3Bh//HE8waNKr4gxO4LTb4gUDaYONHwBiXmCTknYJXgKYNC4+hKk7JXu3zieWdf1tKOag1CXye2
k9HCD7kWzkQB1BzjsvijQod4DGAWiPDQl5XmRphUjBYir+fisTTAh2Ruf1IWIwgiKNrCeQN5oSai
BJvCqrfGIK1nYPiDqcFgsxfLYMa7tyJRzXBzRotjLjcLLWIxgHr1cdZb3r5nKBwf7GAX4qttEqqC
bQFCKO5KtmYQ3dGxu2vvbfIYj+/rto/qal7KDWxEhZAeaXnoG/xwa3vh/SWRfWnAd6pd27C0IiLb
RazVadYD81BdCbocLzK7EF9K9cIDx3R/wHp9QI3Fw/j6c4/MnAlbs62XPYywWqXvOJWvzv1Tbjp0
exPFRUt4U+7dd25Qvr6WWRvIrjvSgNaL4idk6eEnBk0CROcgX6jKmu/3oE+uLS5ZqntH3UqVAHZ8
SW/u1NKAK/lesb9KGOluP1XPbwLlckSCaZd1Ui6EEco6O9ndb6cPihX+v7mn1jZdpDUkc1iw1yhR
o4dATAqB0GOdYuXfLTvsxvtHKyWQj+zjnabrHRJ7KeAnTMVc3zi7ufdBi0QgFSawgsMz9KlfckV/
bo/Pwxm/QSa3ErD7ueHEruHxoijKcgnfiddkoE6eHE6okhQN9wn2/nOVvLUkPm4CERCjNbXYFX4d
Y/HIplqoc16+GQZvXE8Cj7keqNa4PjAk8NiAaU4MU26Ybw8V5n8REZ9zCYK0XN5mHiKij6IINZpe
fyZGIq4Alo0jPd0vteEm33ktFQMYi0ZMn40vqbjIyNOgn3lpERt5XgIbAmsDeoSy7fAOpQcS07oU
2a3XrfiBULYnMlfEkrGCwtJvpitVGn3FhPv+AE+vkgjtW8BMLkf8cL0xkvrMnLrAFX3SXdpu4+WH
bnGuURB8xYLdP9//PczuQe3eZTlg4pQnqx56z2OjSMY+by5qh0u4AMFokc55OL9hDwk2/P9o97ga
SQ3soG0a8F5HrVNjTQO8Meuz4kJX7JohkD01EmYbt7PTljIIxQ3M8obMwl4AdSakZwQ9hUHlvaSq
vR+ti1Lw0wOznfZwIHToh2NHR2ta6UXXDOn7fpLeK/jtzGEEPtmrSCjVo/vFmvzDXgZDuCQeEpUW
uLzzA0rzFQfF/i5QqDFWBwyK/PC5pMjngEU/SIv01lHPGGUE6OEtRZ6hD8GHmmGJVeDn27s+E6WW
hq9jTwjoKYrjyPNrdan/U4gZt0gZR+txZJKjMSCBZ3yoswJVjsXW43owe9gAcAHg+irj9yAAHIZu
PwTEh+GkxN3dcCpjt1uRurPUKE5k+oeU9RK8nlfrQJr7qA8QiS36DaenZCdAr0c0/r+Tq2V+K5+5
nML52RrxNK1eJILI++tweJ3bETEx3EHly35Nan6KU/Pl/xydIKVGyWBxuowzEwERby+ETk586++A
IMBzLtEAnYNSqMeIgot0KBZbhPLDfRnpqAyrLi0XuJXOUpBWTQ2RSJpnqmYYvV0aEZPrZDg7oNk1
n3fHQOkPENgeGxdn7dp/kp/k8MsddtnNrLlrLm9DiJwas3BQ6Gj6BZ1bmzdT2swU10nuIYF9QROU
psaHgrTz3o6Zzd+xsnklZk4A031qm77s8IIzbwe3WdWhl2KVT7OCWwRXUFzi8MieAJcfUzLnACd5
8hDFLjw9upR/NKL/myHiYDPx43MukP43qoXCppCloO6odPallxrWn6FHRr3HPDoAPuiNDVXb3RhS
+kGCCvm6Y7/PFRCOwlWTFXtn7NXmS0z46J9djGLE79crDICRKkebzx0h9bSaNbfm7WqUejW9CM7q
Jw568Xz47QafbmSzHw9ELGK+LszIRaWpDYqG0RZn9VR5QISSyP6etiXgN2GfAusM8etEzYsdOXI+
NFNDZQ23XhZMbtNKCtAR4Ayp6pIgfn8JnYLFUGE5Uto9Mx2Gm1wtZTAUDbARGm/jRfgUqDstCG5O
CKHD7VKa6EHYopnMOIJeDX5UKbKlNaAh0ymUa9jtvDtUJqfb8OuJk+nv4ZlscvBfIYsCd4U/n5IY
GblAXe/2lGckzLSeAYE7+ShOgmDRLyI7AH0puBXXSQOeuynuxz4fORqVvj5Hx4BCZf8a+f8UH7/Z
lhnHMqX7soMuRVhodjFmAnBSEuBVeydwfUL0DTL6YQJcIinK7X4QqS2RvQ+BlbBf6l4oFw7fi7sw
7grmTKEk0wYXO+LqaGXVtS7M5OCHITeUEz2pkC3/FZ42mqJajEbuVsziaGV3OqPiMOwvND16ZN3M
J8dbKq/3Wr47uACNHoCRN71TXnFNIea65+4Y0TS9VURyeitJjjnqnnAWaHnVVCS5MzMZH82idi4e
gQdNXOLugeAB5VWEEVF4UgeUWI8TMQEECWIGJMOKrvw4kvr/k73atPULqv3NlZvqK6BOsU71sVVm
5gBEvw1cJnRzFQNW13xQcNuGIBTyT4IE4OTPDGwg5b+8Ba5PwJcyIN/UQ/x0yc2v81520Gq0WmS8
Ylb0xt2lacEs1pgtcIucI4nJM0N4/kOSqokA3ymuQ0GXmS7yoLC7Nu1/pOXd4ypuuqWalaT3itcT
cgutKFuQQS9DvRY+oCobYU9E1deVedxIQy3MvWKKfmhYg2JdfFDa+aTA/x+X8OVCC52EcLzMxJxH
rwkupCTJizbLo8TCF3sAoavjRcOlELBcsypUsi6mgDUCASHrCuN46lO/SfeSuBCY3XsxQl0PFoEM
g+5p2gLzQesdkds2r+nJnOt/bP7n6ssH2wIWH5ls5crfztJGDeVRLjfd0koDShHKP5zfnyNUh4ek
ZDF6zK254RppPlnCR9WclZvdZhqVwUThSQpPwxVqR0HgR6YPki56UZO0op6ZwK39wAWknQA7zrdL
N0/QYtb3WxfXK+wmdpqp+cOnLbY5mN23I0ZdPHAjAPbowDDtLgN70TOrYWrt6jx+B5jyO7XC9lPQ
K6d/kX33qcRtTsrCJrLAGftSZ79dHzQug/YiKcJxsn/645R8EpITSkucjuY7b8wFMRKe/HvmywhD
cVFjBNYZHUy0PzSJc4DXwTENIq3jrh8xwhk48JzEQCfEdC9qk8S8toZMl4T31EHXRFhIqOjb33vY
XlL/fjnSGK5NlwnkXzlbvOlz1dYp/rBA8XLnpgcE3Jh8NInzGGF8UcqGjxlotmejI1hKtsVBZpvn
uB8rCUW/fITPPIdU2U0KaYDkaXaukj/+9ogxnLdTIwezFI07PtzJrHWbKri6MvWPZY994n0ab5H9
o388QdWgxqAvqZU+30R4nWlBFjwnZ/Q4RyG2wxu8V5+1yHskRt49Iy7yEpThEuZAGTGxw8aLfClG
NqOdG3sSQxwzlBVQWd3TVKO1iveOqTDxsuorRNBt0dGX8wXek8lVJKDKwDpBjydatZg8ayzJvqTb
VKNpWK1YsfVeBGW0RDbwR+0d0mJLiT2X87/c4/5ZoBzFpAHtKZmU7Yqupl6HqYwLPG6ls5nl3rxS
caNm0UTl0BH2IWv+Q71pFMGimL/Cb3txfmIHTuuUMCWEtIlEy92wGFy7xbyT5jId7lm4CUuyPHbT
2k3i78/mgImef3902DMDvsO/N99lX5Ahr1Gpjh7KxM1ZH/93/St04XW0qFFkN8nvNG1c9Khk4NGP
042D5rmlw4IwXMeq32EepegO07bCR1krPVJedkUgsmNOX3wZZxFIGHr7ilrOvhReflD345GnDBEq
2ag34bRWxQreuGyABGflXQL4IX5w7kaAO7XaBF7hag0ZrtVkL37yxtX4SzAu63jr9qvZLZhFiRT3
AX+p8qndt6LRWl+mquyhgmMUlQudi7TXSdujE3kKjBIwG60GbyDQBotTIe/SjT6Nxa0CFIa6j82I
A+9FNe3kWb8BnNByVYOcjM1X3stHbwt+4vyvdYx95YSWxcFgFR9y+ZRTimjnzjIGd7pJgsTjuJmt
ZpL7K/+DOK5Idn+51/Q1D16Gr3v28tGFfK4LOTutwzTB4X6doELT07ty1vNMKk3rEoHemiRIlaTr
sCMjR8qihsDiCX24YWqlogSLujiDe8bfKITDBqh4rsPd0AR7y4c345ThDxzaf/QcQjmhOliaGojB
nvOtMQ6lbL89SzL0101XkOk4l9acbuk1YDRZeSVpI9nloLOr5HpBLAUi4xyn5yVzJdQ5jhGDDkAZ
wTG6fvN2GelK2v8kqAok59ID/zl73ZJViXTE/A12/4UtVQHXG99gKJQr2QHECb8unN/TPvj91sP3
PW5k03Z97OQgD3ShpXGY4cdYdIOKeVy6ViQM01jPl/PPin9jW7VCXhlUvqm9Ub78/Hn2LUaA7NrP
IGQCJD5zgFO/nngItQi87xLEGJ4C2FMG+CMV5R2WVfbEmGu/2x50x0txCvhVnsHchdDxIPc2kPXa
h8vXs3/L8GVCgbSgAM5rSQMgIF0jbLLbP42hnpv/0SLc0nVZU6Or7NRrYCnPkM4/ccAkkKG6tqNN
e0vf33WqpZzINFzpYMF1yRW6pEjYIv8IUU3OPgT3oEC1irndlu1x/+TcuENEz8IY9O87smrt4E8v
kf4MP/u/dGuP5hoBDyFJDtzG2uHIqp70wbZRA7mRJY0hZG5y2d7a0JlrpuFcOmXrTozhuabPVpUT
N0Ik2LFO8kgi2pq1FiA8ihGuUp6555pRDCSvtTBGpZjuAJj68MRkBqQQCplczsNLaitH4Y5VnBgK
BIN8TjnOANu2pdW6+LSYRAcXO2N6F6KQ9X7pLnjinBLc/X1AqoidrVoX1AYDx/BEWTxMeQnBle4X
Kx6ILfVZN+Nk1CR+L2cyuFYIhVECxKWtSblq8Pg3swzi4o+Bo7Yy7kEFvxsN6fLAao3uLPkj88D+
Gg/qfpjvZJEm00Kb+gUQXWFkiZbP4GkokE0hjivTLQyXsUdajKvNXmEMpskps4J/ht/VA6MPXhDt
CelIjEHJb6HIuhDZqZW09oDcYv1A/KZ/0EEWYoghDlo9BgTl6FJhkSlAr5dz7Q9O2UbZbsZZshmB
HcGmIvqoY+O15hDUPGfVVnDyGI8QU5SpKYItKyu/31jq9h2cCw1frJp6LYEjCiqTc9dyqMjjOJye
HHJmIl/hCamiEAUqpo87OPgW/+GImGS1WXdaDjM+F85sSBsS7zghcS3cr2i8XXKDwHXKYkFN2rOM
jPmlbL090Hiz8afnB43U4i8jcII0igIZdIomNlDsJXjuX2J1HVXIUGVwqKbyI6oyCiaV4DKI0GXj
BX0yH2LdvGZ+cfrJjTuLkVuVgn4obXuFoiloXeFCB4+NX9b0Au7RSI3CBf1l6yy1kxguRgfmL6ef
FTidzVcmGR7nFABGq8LNbi1Yl53Y7t1vuhwH294Dtiho1B1ELMxflUtWxb/f+wmsTL+3JfADWxWf
QeaECxdHTdf3juPkFfdZxFSrw+sEM9MEEp5SksDwDqYGER3ZPpSTP9JXE9BtN+WESQRjsG3F6DRk
+9c4Vn5ySA4FU0f8ti6aJjYE/pGm8jaEDcEZ/6DKIITS6JsDelZE23iIoKDUQpZ1TtZVrR5dFRbM
NCdhEKJ8+ixWx2A2ZFWIs2pER806cwccSgu2iqGyz/TNsXApENPM37WeDBjAns0xLkaRS0MOhJjm
Ys+bX0iXmeDKNgj34Q1Bup+wl6+zHNcDO+Bu609pz5wODiS/dpCllDdjPkGesUxOGZLIJUUlz2ub
IAUh/cboyO0QCMSWuWW0hpz08sq2oSofXAiSILBhqtZtfjmdVx31Llr36QyA2KRVYRy30MAzc3HW
B4fZQ8zL91vDcCt8/eFJLSQn9D4FafB6uEgW1KhkihRJIGYmVSH42lhU/b+8qIwtrUpV4p60/FOU
AYkbrZGjhyElChvM34uE0BctKFHn/QGEIeA5P6TmvFE51qjqaCuNoJAl/yDDWz9SwP8k+OVeCsld
StMs01LTa3BG7CQ3m7f/mLdLNyK7X49+XUCLlW+Zaq6HCwv2gA/x5htD5MmYa8nNQJnXeczIXxNk
j38bu9UBx/z6ngQdS8PRWt37Dpd1XXTd8fyJ/m5eiEORa4uohNk1M6c8xrmIEBWSbaH0MqiAfoMg
5jzcRIF8N3mUm7xTKK4LXu1KhUoh43iYO2myfuq19QWdfu8aGtLRq4kMaIhqoDT8cfuV6ZsP1Elb
AILGOMNx1SALWsbCdb5Tz7YhiSdOWaKSDMstQtR2WjDSLfs/M4wcWrRRzUugwPN1RCPoSAwVTWF4
UDRsxlLdfOq9LNVbRe6Yp8vk2boT6rW7E6eQB0kT/L9aq2SbbevmBDL42cXpRHTnMQEaGCTDeSWS
fcukdCEjgBv36GKFwZui6wHJyIhxzcczZBgXJzQaa89kXgpHmVQ/M/2kcoV4gxVi1reyRRm1DY4N
Ovnv1MD0UBM6srFXJ6zzDBiot/QbJP404LxSXDmnW8+tHK2OkO+m/UFGpsEuZ9xZonkyGqr7SXDT
96OtZlq/e47yUWZv45pQAZQY+XRcjtwsYUlG151c5Pi5+/dyYwf6sG7PlOuI3d4LZJ9ZXTzh4/+6
fKA/51Hj1V+a3swiNlGmttq/PSFKIuwd+kXibRl8C+v71+BU5IRwavid6MJP5DUko0lRiGUIYfuY
nagwxvxDbbspaLTkmpriM3La/7Q9LP12OJOeSgw0P39i79ToWeuz3YLo7t/BEXZ4usOF/wyZoutI
iuEPkmx3M2wBt6/SGOFIkQ3eArWk4odbfxwHX8EQcwswDVfMBl1qeYWdaOj860V2Aa9DPMFunK4B
xYnthkWSbIFyf3+wLywS/d0cvXvg4WkTR6wUB7nqO44T4Yqufw1dJ5Qp1+7MCFPM6w+RuHspuKYL
BLrwby99hJrDSBr3ga8oOYeVwv1aw9PdKg7qTLJ1Oie8xLxfpdDUhNyxwe9xh4mi8przrX0st4km
ETQq5jGtx66FiryiSNegHinSS72GItGRD/XLqcuhOfV8K+3n4ASkISvsYBQIK0nEY3Zn2OW+dr+U
omvVNoe7LIek2lMRfn+cl1Hx3RFbiavJqXFxNyI2H7gfM43GbVAewYVpyVfcuSEtfvyvPeBChmDG
GgeBnugDyE4nt7Kw1jNENel4Nu3gTb4i0rEeLNROQu/kHyrYqHg94rYeYlXNC35CPssm353bLXwu
wbVHLFrLv1gu5iQDKI478J4pc8F/+8VH2tQdcW37WNeH9Uce4wwEItADpn2bja6zTF9gI4LqgtQX
AbZRc6vk69JIn+9AL95NtzFcU29QvcSSGohHSjefCg1CbiL27edzCb0R26vELK/s61nAgfIkH3Qr
ICdLMwSiCs6pPM/DT4QhalLzufVIWD+gn3TGfiH6IlCfKaHKn38GmlfqAc+Ytl9+ePkCo5uFEQP/
GdshNOy/x7Lyq2zBiCE0UC7jKhT5SGMujLWR6Nf80Hs77qqDjnRo0ctKC9vORPQS3Sg79QLirNip
PKRXpm6Kig8f098Hpd1sv7EPXhCr3eagfvAb5AbMzCzXxrP7XwLX1efwVW8qVB27okH/WIxyiIGn
9JF2mvwwbcADmxX91XbITgahmmyaNvfwIwH9TH/OvogfzOo6NFOlIPxzvJPrDfWhro/yynKCqPGs
KLyf3AYHiNOhkvGCtiVWIY5FqVMYNpLRYor950rOG5F51ldygGSpRTLTuf07ZXa4nNHy9x16tA7r
baxaQCooRxEcClJpTHq4eA2LVB90PWqLcLarbujcy3LYfnSwvhjjPfNwwTKSsCkp8uwpXOjE6CrW
4coMEGsL9ccza6blRp2dMswMthzvfgbvpLjs2v5cl7f06hvUQvub3+UwRkV6pHJgptf181Myyxo4
nMUDBegvW9oNMetQvLc5UKYZs6DHaEbuC2ScumLWB4+udfJv7qPLCI44IPW0k/Iiy7HLteggx4Ir
rFsBMEy44AvmvOPulxfIMgw60jnj3QB8zKY46nD2ZpA152W2/C8IvTUVNsr4fLKxb/mL1HeMhfPx
XezjffbV9erfBXEyI79vqSMfy+fPEOPGKm0VdLQHoh62vVDtAWBWGJN9U4RUH4wsoqdoymAHhhML
AxeYHfjyd10Q5f+OBAluEJAyFED0osjKfmsR/ej3sFs1tiT+vPNFWDsnY9dz5LQMtRhnfXZ9CgiC
9QqwIc83Zrfvj0bSUi9lt0alvHWqJc5yUz/lhtEwi2qwpmiDj/c5cB33UayRPxTQX77rOEjJS55Z
jz8ozX8aVsgDC2uwffOCVuqW2i2x610AY9DE4wBQJvxg2wuRAiPAeM3gDXEdfyjlIR6kQdwBONND
Gbwpc+DDTN1mqBGev4WxFLWvLLdwOP/k+HVsquQn/XpbBlz5inX30ANGqTsd2ERZ5eP5s9E5fHJC
Byy04P64m5R/UN/tk8c6XFqXMkbvI8qnWFyfy7bE71KQ917ft1OVLEdFVA7yFMkxgHA+zp/XQ8fX
QQDdS47NAuPnTz0sKPwCJ/HvvhpI1DriceyQ2Lt0cV3Gb2kTRnoq5takBYPAuKBPiFNsHEJ5hbRr
S4k3zslMxo7sN8YH6dZ4ASn1vSxjLPkkHCq3mvxx2Fx5DRgqXn8CZ7S2mzQWscsfMUppRcnfaETH
f+KJqjsG54kveUCPwe22IAwQJbYqNdJiPJHzo10cKqSxS3RKwvRGB4IOeTaSbwbWgK2tKZZ7e2Ip
4YY5xBA0rLlbnIXuxqjI6da5BEU2hIhIFu6Ig8IY4fzZ7zdboe5qgTRPWTJdeOPEOk6gzMNIOFd3
lIOscNfDGQxdsqEaNoOm4SIaLryunx0bBYdYSS8xOWL9MoGSfEUh+2lBCj/6cA8BVCd5XfjJfBZ9
lk2Y7YYy4Q8R4KoxrM8fY3k9CeFWVaZqSLK1eFROc6BD6ykisiAD+9MtTO6UDheLK6kkAEUb6RnR
T1Q/9BStcyc228cqFL0INNcgIa13ut+zxeYmLki1monEK8hjPrTbbROWYSll3sudYkfAQYFn+VYy
QN2ijMBra6V0H8/zkvzTXTY8Xz/KSNqBJffv0l9GEzSDGWk55WA6Xzzv/gEeCKSCKblQHCeKbiEr
zIr+/7t/AqMgQZNEvneLb4rQ3Tlm+WCte5T6iIy19BeOdik5FauO0Ey4LwLwinQ8SESetd9nX+1D
QaOHpDn1UHoAuyxAihlguWAvnz8egDVEst0uvtvdxcbQOU0XnF1wH1XOjqHuHORAU3BfutrmfLWh
1HCrLweAjn1jVSAFtISLxfA7zzBkpVYUDcIAIOn5FlhlRyNa2+H9vBBm/8NuHGUzmYwFxoLctntk
AiD5dMdjsnlpVdxSGHVWLVoNUhgBHKH6MhpNagP7sCP8/spzdxH/HLuqvUQPFU5YHC88jW75JZej
9f+2WpKOcqayTFUR7ljOqtaPESLz6HNEpiJCviKQL9y5iZo5lmYMxT2jDtkoQy8chvFtqGC0rScY
b7WkOBNJqW+6EnYoucIy355nKMEHv2qr/hPMOkChB/lSPnOKVNH3lVba2YDkMMUDFdESAX28K4cu
cb3Hy3g03vWpCjqpQUVmH4kFFfTnQ6umoWtMUIIAVrbpDXFKQaOu9BVwoWCOOyzIX2KzWMdViY4o
aodv1sB57BRFHNQlguNhpKb7XFU3bnu6MZ2pX+Uxvy3OwkMtlLeg1zwwm0Ck/QyUHSLzHlBNDYhm
MvBxFNJ1uFt8ZBGhN5lqKulhhJ+PaPe6AgJMa+IefLq2FoQw4JkUx5nCP63FGBdYtWq5izsn/iaP
p8i54hLTLYtel0FonL4XKcYaXTYhaHVL/AD9VJuPO2XFxa9Q2QWWhuQ4ITOPYeoQFlgwOeHwToHz
7Keuv99oawzpk2UuuDdCqo/cDHd+lrIX9pBdnJjA7G7labw/rowNwwkV4QD7O+Q3bcMorDU91o7p
zKxkw3Zzmgyzv9GKSLT7O8GyGaG1rQ4bcppYkRPDhulvwU5g9uZiZEpq8w/avx1DmDb8bPADUBfY
7IqWBYHd7in+F3CvYL9YPhd8rdlKdM27Jr3hm3cpduydE3MiMYW8g+r5d77owyT+d6mvZXevznSL
Xfze4ppvBhlhoFnl5orwNGkSY4J6l7OiPSkYKincIxuOVpcUryCI+ofMYk9QSnk4yXtZRWQgm5IC
EKrf02CNW1GKoQqg8isDmTbPK+uKRCfV8L0N1gpaog5zMzVuIKW73e5PYg6TZfhfAxzai6kd+nt0
SBlHiroXBMpfhQPcI7eBAmF3XW/Bj06K8TJheumB8TOZLEDWuKAzWznsq85zojIkkB0QAS/yXgmr
jyUKqOrVjoykPAlo9uA9JFRlmRf4bKKiu0VsSB/z23KXzR4807MtSuifVioLTi0ZfdOp4lLr1iuJ
mVMdUHHyehm+aWVNrFRfs+k+XBPcamBqdSpRgSUuYr03c9Oy2Yk8WHqV+Fh+c4YO4xv3DF0Nl8Cv
HkI6vl2Rv/lac5+fUtCnV2UUX0qEEDf/PvJYF3hNOBP6nPSHwx34NslcUl101X8g0HTEOwA2LzHJ
ASJxflcchQPeMcjeuF8iXBngicMA+LRpwvp1IlkmWKk99AKmIHOo1u5ooruxwU7VsLBOxpGTxkbk
HorqqudN40Ga50mZxUTAQWj6/O+7LPqhjgYC/z3bfsaC7+1sZ3979MBH56cv/i5RtIE+Mw5yqyfi
gSmDFQH/5kS/bAV0A+OS4yse4ODXYp4HZxHR+KE3CvjAuHfzlUWq9j/NA3rp0+AjYzr3enuXHqcx
YbJi16358F2CiVlV83CtfZtwamlIev/hgUGB5+9FOyOvcX9Tvk6sfG+D5yefGqjpgjY1onFRm1t/
JjsE4TK9l9P8zKChYZdORufp8CsSVWN9iszSSm7gGhqlOXHW8Xc7MAEVsz7Jsm+qfI6017A+fh9e
P6oPlH6C2Syr5oSJNJonLzNfEdjx2tHPrkWQyMK4zkQ5pdf4pc6p8tipOEE8K071S98q1lwUtJIm
fKUFHrBCaWqe7GnUaHEKFmQTZ77hEpCEGAzk14oUO7oUzIBISgT1RbVXm6JSBEjC6cf/ccUgGtvl
7z1fN5/pYBJqt2py3ImVtwZHYMSuDwkJmeHzc+rReMUsJuir2x9hNBcdZjeMWsyWzaIwMzz8MC6q
Q+vfO3kpsF22XwUGCjOrIXytsrYtG8PCwfVN2rs4xJm+EXe0AaevDoKGPAvcHPmw4ZHi7tL0VXr0
3rSt/zRkOuWJGRZSo4LvLO90DXe4JTL0jXk0/sGT6k++m4pNXarFuGw4qKb9PWZBj5DwH9PIg2k+
0JebjXl5XdN/Z3wkZyIh27beVHMGqH1WXRTU6E3Ju4V5wbVFoIo/xWYbkaSm/xvYLgMy/thBSDW9
wMzMOKRQS0CY0fruzM2/6MTpRaiku2PSUpeiC94CwYeHwu6km8djZ+FLB6ZfafRg3LrOXznPETHr
vYmZlzzaImso7Ffi3n7olWvRiwTIOxEATLGEvjvKi0R8GZ9FeZlYcV7z9S+jfPw2jDqMl0D/eZ9i
Ois/9An/dbOvx/AqSHA7L7qOwOjHDJTxlwZCdfPiDUSheyJU0ThxVb3Z0wZHJ6RjnagG41kSe7Wt
hOGijoRPIe0nzF6SG6r5982tpBwpFgCm+zIdB3GiKHsbkTydqhPGKvSoaJlaOh3hb/mQrDl2aIAL
B4BXBRDkC03rhz9jOsNIM9YzRmzwEt7hmT8YHasILQnjUEbVphIyjoxFGZ1Iufkz/VwJfrNqQssU
41kGg+BzUKcjuganAqnPb9RyNKUoraHuVCwmDykYeJYlt0cJv2dWiCFdXaJHMr8f2jX4fOo3pL/5
PLW+PyYhdA8kyk/LtMZ1qjxFjhG9kOKoPxbJmLaHYoWu6tC7H4et0JByEXIV4t6Gj6btrZQactin
q41b4pldCp5JSqxhx+wFdW89GI7/5ZtlZcGKBD5+2Zq3rLfIvpK5d7GXYFkEHJfQwKtGrl6i0kHU
+SmOJm0whtKXNVYvA+aPHSthXWAjOsqU5hFEUIZv1tjA2hX7xjf02WpC0weHM2z3L8jQ7ivSdSZM
890Ilvji0ND9oBdk57gycm+Fok0O6rg8TKvqXSLmcZNGnfCc/SYTRzh1gJC7UVi997wTPFAOTlHm
SR2DtDaf/bV9VSKf9Q/n7sTM20JUJpAbMPQbmrSjt9xRvCEBJC2rTRf7/tuIjin2OQbElI6KQCtx
x+F4FNZV7jzC7Zojfklt0ddtYBE3VfdvsGMFFi6bkyBx/wYjYwK9U1HAEX059fB0eCXHwwIYUQzL
j4eBx21BkyHv+2u1tJgYkeqAaHSmfRNYxyFE0JlUXAKnsIM8+EjiWX4GDMqUd5V2cbVlPxNC8/Hc
pJe5JKmOdwz/TwgBwA8OO4OwwV9ihZqjSKIgbU2yHpUrZ0spL4V1l+8dxwpY13X8kf70i1KbfZFD
gtiisfapBNRIZIIOojW3IQFc8T2rpnNZ4b6oJuKz3+9n6HC7zBY0wxwDXfVZ6F0JIChg3b5VhBoO
gzk9ayZCU2k5ij+2m5DjiceakF6P2Sv7uGjtl5wBfJ4/TDCB15fLcPD24WYBofdGRpRaKvQsXP7g
CfEveuFU4fFlVewGQgfFLDedoViFdqnhzMzg5daFyVmKmq8eNgJx+npjGjYbSNyOFiSbcfom9Oeb
TrR5BuC6G3UByEdNvaaYoGoL/yAmS2vdOyQqJ0aGJ491kkHRj3Brd8IXJ/cxp27/OxZhfG3y2dVS
8FUaStLfXPfLSOcYkRno9fNPe2tzKM9zgWXNLrN/iNGEHfZ4SujXjhnQU4rpfNVRay9mil5JhOXS
y0wLd13J/8Q5zFTIaej/HpPG8JLEl5ayIljl2GuLGCiNSmve+9CVAtGVqlrRD/Vw6weblFoACAti
j8oMd74mM9GzCsoXyjI9gKPVYvdWkEjPntwO1C95kZdCodLaOnEa1zkhOmzGE9MMZgHNd0m0Nrnj
dhD5cdwXLMeApLzp3ieMumUcY26bayKbsNlaIrTxtdgQ402BLyNFbVleICzHXBQ0bFRjNIAYZaBs
FxYdxq/cMKT986TQ1TumCpVZyTZfE/q1cLH4a8pp0rJoFkrCrxDkJ3R/AaThGW26fKwcij4RaTNq
FaKfsdH61DrlHz8n1+ygNd/oARiYLq9/OGXHx2OxyK4JrwqYsUmYIYyluGjI7RbQqIQLudCNSgXF
wG86DK0qbpD264/mExf10+D6exIKBJxsCfldrcHIEnENM1rRcvdioq29F4UQy13WUs5F3ka7h3LB
nM7IBneTocg48ugmTbia5+3wDXao7qC0kfXF0YfHgddyotmhlyYjAT1kbNmGPqiIYPUaQ+wwzroY
+IrrXhtu+sF24Yf2RUrsuEES1z16D2YsahCAfxti70rGpq8du+ZzvTDVtNefiTCJx53ZDYghUn0a
Ab7HCwM7vYqz9phr9CCuvpxiDZb/Vb9GBjmF52eh5StjKqD3j6H0jqF0K55XeZRmTU1qh/BzmSzI
q9thNXGmo+9aK6hRwP5+qCTYHyNFVQVdfKvgBDnuFwDBzDBNSalmpppGK0HHE7nBnqigI0lYGRXF
HpMwQ5PcGND5T+ZqoFqmL7vAnGv0/g3knW++/DlGq9/5ouG3Cxm3ZFjjOAoF16upuLqU9jmcZGka
6qqkXLFGiaaL/o5ZNNZ3kxKQsW5Y7graBntNjG0KRRTap1lICjGY9ITs9n3Ge1henpOGYqSf4ZlK
D2Xt1kAXWaUFcRV2pQfLnVt/xQWZL+dgFBuXhVTkT1FV9EhcVDQlymxvW09KsvPW2e9IF63G3Uox
qLcbN3t8c/PaKoOqIG8OBeV6WQqXT3Rc+u0qKKhZUHLTZKX4rYO4hPKNDkCjtZzGGtS62/eyDwBW
8mOwNJPesD+inN2MA/nlJHFrEcyblkXhiLA35OWEw7vSwHe+1wHaGwwVpCROB7MrWEy6d83QyaJr
KQ9uRgDllLQwotgR3zLtFUi2w717mRZDfjlg+/jVHqpGK+AVQ5m1jg4nrTQq3d7Ajz8cAd3tLc9s
IHucMljV1nmhaAJOmdj8CUOp0xtE9HH5WXa+6ARtOPgfOGNFix5F0N3AtHycrL0eZ7Fnc7j7jfGy
kROBwO2YPwZSFddnCbmr7zmAy1leRVGsSoRSOt7yTzenlf7u4PCurvkww4tjvSYx6Kri5/1/G52+
/QtO7+BPDI6oMW6cPKzagoqUM7cE13akpONywFCVDijzn1j2VqCKdVgs7mT9eSwDneqmxVWU3vjh
J1o8jUvoeVPDOyV/nOVOJyIvlazEf2nXsetdk9KfdiyU5FCRSMI9ZPoyb5JEDlqn+rNg/Wf5pT0v
wfPw9rTdWr/kStNIh02dCixy6PJCbbdOVfQLtGJAxMyHI+SNhnomIjIvXfVWLSrEjenfaszFkvHY
iEWQ7s2RBluW/8KD23i13VHCRUdtEilQFqNnm7gdTdUNadoHwNy6IMEJn8YkJ1wT2uEODxu4kkVe
JjZuA1A4Acet9mV4e6Z6aE3Vm1eUIyklPE7c/BonVxlbIH80Bst9op+qEgBHamHeFtSHbzH1FuUE
KzwACK8dWKb827yb44JO6spjuHzqmmJolGZt2edKx/kqQhoCLd+tdWibq2zAgd/Wdy7YAIW/GACq
X0QjAYPiuAXGQaAmrwf6bRdN6c8k4QrI9oNaP6zqbpYR7gZhaEGTpeFBfblqc8Vl5nI2jH+ekddN
BkmR+xg5+ZLuP94Tj9d6QHh8IFRfXTCpm2J30SVfqcgMqExt5/hpbxyevC43Zt+rhJRQhVAxzs6I
6UadmFZLg+ZtLPkPmuxq9msC16kn4AIjBUWeCy0rSafsau8O1j7pGLEfDuXoSnTjaIW40sYnsAGo
n2o81MCHMJJMCUZOrPNz0CJdQLdjhjx3Jw8BcGC0N9JFJQaimhB22ybCQlhH0fZfzl2xfDiPLzzF
dVdR0p20V2sFXHwtIDDlXrHd60TaOYE0sDpY4zMsCPX33DeHYEYIjA87VLuJXbEr6sWGSEfLDRx/
lFlwOvnQKBCmsTBGcs5zYDzANU8RgzGp9Xccwik+Eu9xRFg0rrLvHu93XWb1xSqkF+TK9UuT1EyW
MC6xbNKCJrY/5LVNumsqYMaNPqzbwCVrCqiC2dnQuHYfkk+hC0MzqENNYxkbW1bixDJu22SSrgQG
sCaNHJjeqA3nKKZkiWlnWtD+/lR68RsjBo3XAt03hyOrEn4/eh7vrnewC/w4HHTtKpMKQ7yt4HIV
E+zfpawYawKCr7BfthW4jkXKCKkAFi6Ir2AemTWq4STT40sRCzLwHy2REsubbhuv+Ig8jNcV9/p2
Pow1KLpgxAmNmIWYLv7YG6UWWFKxX4F73ICivEsJokPtk4RAeeEuSCrdF4j3bKIsDdWdCvHNjvTZ
euLFk7bm8uH21fGexItDi4CFOJ1RpaWh9XH4TxUOdeH3cMe5IrpSbLzDKFXE5qfUVPIcICvKmEBZ
orvs6/RZXYODmymkUjXyggE/sPjBqVpwrwYVF91nmRP1/py7K1Ka8XmWslujC54p92nWWX4JmNoN
lQYphApgZqUu2ODKBtB3h+sVytRHgq3RWEp2sYZT1Ac4rjrMedtu6Q/yi3oz48L3uZf/KrdfUN6Y
c8p9B0oEFatctX2ythjm4tqLhSwvZ7xJi8Aq7QUDKaPvzsScmjDGoN268uVuedlWPxYLwYZ4wZx5
B4dXBBNzpVupXkcKXxbzWJoCcXmSHwpGaB5azu/vvqv6zo1W7QFWXxR0bQH0vL3Ge5Cf9kejdYdm
0RUhPlu62mksM/4IaaVyQFYUiZz2oWNiOidn+Y9sH8u0McS025NUa0e8UJ1CxkaVH047F8ULC8HB
QDL6C8+Xm45WvG9t0Aqx+y8L7kxiVZIgGczqLHGCkhOvn4j4vhi83/PWaEzlYJqValPUCgU3msz6
L9b8qWCK6OEZRY+k339dLj+ghXB2FC6VbJ4oVI9zoms2a3FFuzpxRXPqF2cWyDsURuPINAlqJaCg
uQC81Q6L8t8nLhf/Zzi9vjWFeECAtUwxDdpssVKZwe1IEngVSW0A1sLrwRfNqMzvZJN9lqQLQ/p7
BP+up3VlvIIecFOaI2E+xyZ+pPAV9Fn/hmKEjNJzMIeh2CxDM32s1L++f/RgXUMJMcV5U6XjXsFd
+H3EtVkP79cjJ4GT6+hPmzvoahaJkxqPGxRhYuVLW/GlFB//gHk6qxbPntt01gmAigGft2vyQd1H
3K8oqtw+o+3wzgK9iEpaJnUtq4wU8d3oxMqCKvyg9J/RA8dkncZiqjFxOOfPhAeW5pql30IUyt0J
EPPtutLsG2ikUWMMT6CmU8HlHljwG/sGvemboOFlWie38lmxKkrXLZHQpi3PV7cE1NbKrasoDxrD
W+QquMfEvGoigWUONwCg0LLYvl1luvPf69g5V3ZoqoYoE0RwRvrVYmq6M7mfVaK6qeOT5F+LsoAH
pWkcU986J4VtfmU/d2grKjFelIRoSn5ZgIfX9HH8M+1pd4B4mTKaw0F4ksDFTJb/qq1sgyK6wy2L
m5TTPlqcXb7LBl2qxc4Ks0u3wsT8xF0iUTKJ2Ht1sgz+dKW4rHY05y1vduxqB+ZPLiEopMwP51tI
FeNG5Jhq4k6b7VRcTSATXDQK0rRTFeVerROCqIgNg9dYvs/WNQq49VmuHVoo6f7zjGyb0Ljft+2I
ZJ+h3uhLtKN6cNz9HUeaROIdhZIcZ4ke1jJvWqTKrlZPnSvcT8TgrB4Ee0VnJsSP4DIUTQc5ppO+
YXFxByW06Y9f9WDHQrVXIDMUhlId19fdOHQr4eKXJx2KM/wr7FFxZzuJV+4NF4iwNe+o+UVO5iMZ
/a+6PIFPrvqEYgV1nM+khFNgESrfZ5x4RULE6N6vbZEe5x/pvBIsjPMUizA4BYCh8GYNSOeDCj44
vUb+Vw3d7Phf1Ac1mkOUTXGsPEMOqX8PZtZF6CKXX26Xpf3yuHPbmV+ybeBkPHHD1err5y2CaLBi
tLDwMyLtqFoZSUJY5P5JMo4WXHpcih27c30Imo+cozYZJihlH/iKDYARl/biK/yigHQpuaFuLzxO
KipspyYXnEhgt9n6n/mpcZ1VG+qYUwaZr7pfJ22T/+QOs7Wzbfn7qGRJ0Wa6VXt6rzENPkr+5tEw
p/2k7HgDpzDC2bJSPJpB4PD+86+zH6wQWvOvtZLVfFXLI6SoEmey170cdnqaKhLwb8z1csbVRcJk
L5N+IpcvK/TXVk8sh2FF2HSQqONvzCGyzNWxgbK4+0RLHxNJRPbOg9/JonxWC1WeNznhnm++8A7F
VgvIpbRL0DvpUQVaCUgWjH95Q2usaWiKnRUPndqmxqNUjAtKDx7q/C8vf0fqjdPD+o4Bx2h54EH6
+3fJiYcv2uQiPeNlSWrEVFF5rq9kd5sXx3E6btEPHCg91tiTBjHc2sZqsjny1qGKEh2gtXMG6Zyd
uhly0istu+FmalJ2eFiYPftWNKh2nr+rrAZPfCLnFRYgecm7XHX8oJsX1c26gD9zftUwAeI5i3VZ
/HTY5A6SkZMPfl5mq3fk14ZBnjUpz/dwmjw8gvP99zOAfT2Lmq308e1WUp4/CSt8zg07iDUQFQJc
yB0baBYY0ZQlFdDi+SN9PFmbj0lFbt4vXYuc+bk+Du7PIwMbzY5tcKeSpP1+Ou7ukPt0btSD4bl6
dt3k5lpC4+DGFGVUK7Z7WHE1L3+jIwEo7N7vEJ0LJws9iRdlSRo5mWhQkyHwbIfCDdQGBuvs4NEJ
yvrrk/7JX/SOSlKc65vwV7JKvnRRjAA7j8cBjd5aCVcUe3geX9054G2dJsJyVe6rxVik7wwdEt9H
7IFB1+8KfM9hMLP7GNPfN8T4gZbhe07aAe9WWh5Y2bDu5Tm57XlzYAvOpD6qFCBDzMO5n9T6YdHc
7+X30gzyo6BirrvTp3RN8J/KBGWi1oFTPHGgKK/WY2+3x2SWQpIRW8dq09rzk24UOcLT0ZNti9Yg
le0qCpO3EEuZJdy4WcMm/YqRwLloOcZH2iMtvXzWDp7eJ2bhsOVgaoxOOvfHt3g6497RvfU8n/4O
ZcNKIIp1hM3dS63B3CaGt0nztyl3/5mWIImP2jzFFiMRzG+TFMjWPMsEQ5DI/deC/ac1wY45DvQb
9aMrYvlyZS/QqsawknP0UJnQIAva7gMHsKQUf4SMlMACnRTFsrxz3SmVq2RDD1pDpoScZmzVU2ZY
wQCKCjfRW5db0qZwLuS8a+7w2hwuwsBxAds8jp/CvjAaz8ArCwN6g4nvM2F2taSQbUtGAm0Immmw
EVyuThY68KWc67fbDaVZYk3U0ChemXXPMFJxFjBcq5PvUsPXC9uDru4tj2PzISaSkTlTsWn4qAFC
1VEypXgazYC8soN1eVOvQ3g7ghhVFxqPCmDk3xDHDtnbOcRrzCdJgSVukLyRtkJCs5Wc9R2oDsxW
zsVtbw1wsjQm3pMdyu9ToUzOs+qXbehtnsY5zO/EAIvGUzrRyhVtGsYUaLIbs2AHADJCzkpPRDFM
uVQLIEkFGYjRvUQ5QLDVVph7aJKm7EXp5bdyBFJpZr6iSbCCIMJ3uCgfJtMsgkU8Fc9M0sv8Wimj
Q6eb1noFVzL7akjWfTwFEc02Ex8m5Ov0aTeZ+JxC68JjdYElkKAV8q7fDGboWPLxKe5v6HH19v04
uFR+dcGmGHHC/5EfDBbXaon+tOE1FzXMd+zlETd8Q3aYakUuI4zUWgopsMTRuo0kBKG/6tKO5Wyg
STt+1dMNqUKWAcGenD8c/+RqCXOYBP7c+UIjA6qDpMW/usXwcjQ2D76rBS83k0yhvGJiX7TQVDZS
w5v+zy52RxjEjeVWHQZ95NJ3kkIsf2ZP9eg9naMxQjHk198kesy/dU/NZKmhNvevDqLL35vCzz/c
7DPenKX5w1z3xV1W9075MqEE3aVc/6mpW0j6TU/jBcGkjkifyQFgiCl0Ie3xU0HfOA27UgNoPHv1
/oj+GQ95uCJ58oBje+/XD2QJRCOmkUihbzV0jmKdQwQOoLllvU1dU2DlychgRVTYXH9TTgENj7kE
6JgCrcziMkU1DLZhJPnLDflihqFtkdqhZrm0UG0MnV68Bq2BdNpGMLFwTIQCs6tLd/26oW80veYu
9iwzQLzizcBYQnY2XNZs0xP/4sjhSVHOTHtFwFEUfTy3+k0JPSr1ywOiPbKQIHFV6sxTqQxCMGnL
4w8fPMwrvfrqlaF7PlL7m3SOv0WZ0erR1Pv9MA8GsQqkm9cqpoirOQrRsanCkY08BQMSmvPzPoiv
B1ly2Jqhi2b+5PHlGpZzSohduNiSyEC73llszCwwWtlqixVszRJl+8psx07csAb5TXbUAHAUl51E
E7V9SP0m8kel4p4Iw0wo2QK40qpTuTbP7TykgLcFN2HEb9ssGJm89D+gEx0DaD9BEExvVifAt0aL
HLO05lBibBxEgxOutjcp7SCrzESFofQcLhPPebj5q29hNDP/VEf6IAOXND22ElqItD0vkeT1peON
Zt6GF/d6L0/lIY3RShrOnCQuQzEMtHRFCOOSaiUCqOPmxJC/rQZcqC6Q/BgUIUup84V6s9XSnpJc
tKEe2k9RWCuVrGKwdRhVs5/Luva/QDMqDMJAt/FzKll+MvbPyttqMP2W8+7bNizSDLyXGqRSHL+W
hGqP1BncVHxsXx3CcuAVPnpTPO/JrZDjTScwPA0MTttShXsXIm2et+oD5mAFqp9DH1KHYdoGC6T1
AluPJ+810vsUdHHxseLg5g3PbBGMZLvWGXEqfOiO4xmI6LgppZFMvX3iD+r1aBsQZoHYq0eUq5nw
uvkIHOXbF4AqxW8aDCdH12Ggg7IbrLvAI0vVYn5fM47KR7QgPrS9Jyty/W82qqXemtHMI0Q18bLY
wExk/n/+lJlSI2PPhBXBZQHFyl/DrwvN3gFzRHLa6S5vPynFXdT+M3u0WewA/RlFYgy/nAeKljTe
WsqI8EELnjY043PhCx9NZkH8wuX1y/n2R9B6m6ioa2N+R4NRlEwYDDtm2HaMtPsovgXikt/f1/Sg
bSbxCDtXYMDx+Y9FQG0LoJcYdSr7DFIPAEnEwEy8L+XG3r2CAZYqVItCdeqgsSHYcZTM7TfDwAgh
KrgcKaVd6YmK8jMXCUImwMnxPLSEFJQRI8Rj457izcj+4cZDTzYWUkzWO4TdPR+Abors+x/cWXbO
+CHpDnaKggBuZM7y+ldxkgiS5b1u/YcyNZilKx/YQ++5kEyAbVkPCaOkE+hqNvg8ILtj0txaoR2i
ffg4WovJmc5h9kPzasq95P5xqZBD5muDJS3yYfCZOfb72pXwEU/+2Xk+Rz2E6ei3UoB36hkU5Zlr
QP7nFABZ2Lw5D5OmeSbMQZVQdg67xs9dSkLPOZXerXQ1qRXKHqr6w+WE8VETQ+S0dyRr/Fmqgati
lKB4KIHpRkD6a/WuQ//yfADDxA1MwYYOH+begs+kY8YKgvnP3l4QrNaiUKGioU71GX3eJuWq6PdG
fcNfQsohHaT+OHGy1DreUXO/EEO6AR9V3ZtEAWPEO6lZ77fCWrmvr9R31UuyGJZgbmVZbqJfIt4z
9yga4OWCOTDvWn4qsKBz49WC8tMciC5q9Es1h1CpakYLp2nZkqr/MgrQ/fiKSjIL4DiFdPFT7ioy
x98/wfOL26u0vBGXM7fif6e7uteeBHmgnsGM+7zIwsQ2ea0t+1xMIqpSL6Ij1/gyNWFGvCFKR7Rd
hJgtguZVgxfjty4zhuvL5uMvq8RbascLoyvxlllEgXv+Q7fz6TfhmdblGOzSBKf11gZ4itTwLxjP
zM1zRh8Stns1TRgAKqGtpf2DWBOBqKoXwLOhJzK48MyXsV8wXx0ILYZaGEjuMvRGHmEh5jOj6r6+
33qSg/n30hMCzBkpGC7/Dfh7PfwzueghC9sDbYFuvJkdRGIkyWESohewR6uzFK8gV4wY4dSeZpaI
71dvA4QBy2fUi5f0hVhwacJlQjlwyfGCxVD302my1qut1Oq/8nG9gvF6TESRJ90Uz0HYov959VjF
Bp8W2WGmLP1X0tQt3oQPg/sqdRgVY9oUfyLehRJKqKbTkegbAB+DMq13DWWTRWCy5QzoRYO5uT2u
dvLXwA+7sVvApZwhJc8qF4LJXVf8WQCl4iXbN+J1Ggzidnkutc2HXletXOnh4TeHVYHr9BhMi68Q
uPVJ/mdB1HevzrtdIzkmvIE+9ogsA3dPhPgLLy2M0SNaKOwIIQWwTwZd/MJbum4g+GmzTmFDjJPr
AF5hHhTaJRaKAlz/E2zsWmnvbHFxk0skFfnT/DI/D1tjOIBeIpKRsBceOcl7sFHcqo1AQckkKAWH
6QJ9nB/Q5C1mZDBoUB2w6wrbRfD9zdiaLTC510HLtAtZ5AC1ksqaVuz7MYnm+a89GgWE/k8EYrvV
CyRhfC8LYITWADrc3ABiL8ZiUBvu2pU8xDTNFWrljkhHQyiqLowsMRoZpKqp0ZL+mqy2hpeHDL7B
8MSw7SLW4BRXGbOLfmaJp552qUjVzKbthdDnEPInBct49i8B911jqTzpJNei49oVlp5Q+wk7jY0X
PveySk0uT91Ch/bhHNqtGa/fS5LH0RdCWcOtUued+nnnqpaOMTx/XDpfLQcZ5i2YDxGrFc4PDhBe
6L9o+QNIxJ7E6LDpymaxdBVI8UxeGHdZdtVXrYKup8dMbQp4wELolGUe44ud2ChuMp9zS/vDZpXO
9DTYZcgBUYVunWMR5O9xduajwYi7MPqD28prXHVJ350sGTQJRkv8Lg+PGJyb9eltzFPE9JuGBvIU
iKgfD64z8u1JoCTpWY4J3H1mXL7UMsr52QPO1Kyw6E0MWuLWKtPQs5YU1sFKK1dzi6+1vKIshKCi
SFnXsUg3dVHZ5YbTlmpW3SUTMLd07QMC+qhgcb1mh/C2SRLbWv2BxxPWVYfLjSZ9FLVKiNKeLKPf
CK3JY4ryhLtmSs9LHGwpWC9xSu2J2hUblnRimIO0IaUs2wwJigMXxJc9K7pWlRCc+7Bb/pbt8pIW
bkI+IwE9ZTcRZX0Ar8N0EoPT4XdlPhJ/Xx7FeL2BB6IDnz2RE9tys1Of3VrG1TaVT2VGzYyKvtgT
PNPqkxGmVgkQUI1P2aAHcl4Kpb6mdmn/IU0nHdO9lRl1/+60ms6U33qMiMI+t8ilhfY15vp9TyUq
tb049ChO8g4M3LaaUfLdiF0I2/NDaH/Vk6wDJzh8+CjrQcnJEao2aq5daUa8XNjNZ1QnwdU0XIPc
w2uQ5T6trr1l+wUJsZhSQgoG/NxgZxvy6ZuS9ry1ZaLTolKcoyxAP6efVcX7IVOSgiGoG4x1Emht
Pdn6oBuy/DZWq5rW6l5xD6iORL94L+7pCmECASNrCBVpQnScLBZoX571HFRrbIzt2RjwQGqMMqD/
pB2GvKeeVRLq9fCRhxZdO3UjkEiWoZAtImBHekG5zD0MLBHOKZwpjbPY91ahRfxGKYM3wEhgcuab
eUUY8Yc0aL/y++rNlLqVrlARShBJYvml36w6AI8T88PMWkNisPYt/AgnfuuKD1Cpt5f/mEYYkMfb
e1dUyaLh3E2qrZ4SDaqfGmdtnHOW0s/rZU69+sDOBy15deFqCsYjxlXvF75SE2fB57MvW73bKF5d
OXq7ppGj+19rY+jBhdL5PPjex1piRZaz7m87LGqoA/Ts5rQQ3Zr1a8Qzm8T7gpAuK8zAh/JoXXrO
AlOSHQw5LKCMUMGaztbez9+LCjHMXGZOXMbgNFtxyF4TFBrKUHD/P9ZSJnDa3SNr9LI8Ojbpg3uG
vCCfP0HcnjqbSxIHAXzZzon+inGfCWfZKxzSP1cr7ksMrcc7CFKfpL626xKZ67G+8K7Er7BWO/a1
L83qQ6t1Qhatu4o6pHHKa3KW0OcmSTFfCEmBpn1uB3ucntqrULPfEY62gtfUjeInN1FhPEExA8NR
U9+yTHJHpvFjeEWPxfSdwWTi6N4rnqVlt3BjJZYpACcSuzPErVuYeF0HQbf0DN/VBxmeAT0+lJHF
ULGkdvx4aKiGkiFBls5Y80vy35N9fKSmpvv4zUh9z0qmeF/oytZ2PxM55csgx9UUiLxwG0vTs3D7
97gXVEE39QfEtGyLcPPAoQ2xF1MQmr9yclpgqNb2u55gHbZ2W4En0wK3GaZ4jmeRWLizM1kEPxor
ZMYmlDJz20s173WcFvr6ZBqZCo8Nn2WP1ZeFFCN3vZscv0xWe9rYgPqTMbnGiNc0pKEUcMkiVMwG
c0yDiNedYssQioEKaokwTWsWjTUPwlIXJGap17z0tLdqVk9UpmGSGEixJvz1DVoC9wvjJZ0FEXcp
PvRde5iQUl+FXiCQCqYa0+Yg5s/OLYt6EqyjAU2qX375QH46JdbictQAORrhk7T9g8XesB4zAQVV
0zhPBVJxzv2cp3UnGDF2ljw56+5KenRNMM6WILwjqAHXJ0z5sAwz+NwCJR/9xz0dPNcutlz0Frqe
xYs/VPdE/fzGkFYJ6FLcsUc18GjzDl4fo3qP1rohPNLDhIe800igNLdZAGj6dGBdM1g5vJJi/iRP
CH8NAza5tB2gZfWWie2+QOyKayntwFkxFXNplGKiG+4Bj08WX4/GChNra54uuzrl1b5mECNii15P
Qk38/5fG6/d9FkpORsnfDlaBDGTrTyZmBIDRazitKJRi3hIZSj2E73S297AuUDWnni8uol/TGZt+
shNfX2D++Asae5zybTCTeDe4apCk1RDAZnzAiPbYDPPlEG2+DRHGWQk2NYwOszF5JAkeJ4DvBdx2
GnCnZdADZBUf1jrbH85LhYj5b0jjIwx2WL/7s/FVeoQd/Yay1ParuYHq40fgcUzAphmN0J2kLm48
pFV45W9zGynyGhfBCqy1KDPrFYFh7oz7PMKTYpu56xP9DYEpKmmJ8G+cZx4LJ9z8JeUQTfo7X35N
0b8N1bFeWMq9KyGe3hNGa3+JTZFEXG3lNcfp2ivE9oa4/zN8dgfkhXXljk9CyyOxtLVvmxTo0UYT
B9SkfCt+yFwprAvzk25URIvvVc1QRIvbps4Vox3OwLVBr5tVukW7OKHQx3Hi2qZ28a/KGre/1yS6
MYYQVrn/86q9uuz4G3vN61tizsSHGqwZEHyw8Z/VgWHDf3WpeExuVPaEBNID+t8Uigy1PLMr/k8I
0GJyyfPAV84clefLey5045G/4/o13wzConyE1Wtvf2+FeKbMuDDbOSTe5ncufaEJ1yYV0pWuXMBl
RP7S9tsbVx83yvTLCjsnoEPPhrL0or2hVW1Ra4aAsvnvW/AE1GGFG3TFfmuYlrwUY9AvxlQzyYrC
QfVlJmAPAkiFuSKmCp12am2kHRqPxIoAqacxd1xvEpu4IMw8fbx7h4Y+2J/CGWbRS4XE2JphckuZ
iQDk/cb3Pl9XKDGLJwcMchsKQHsfVRQdGS61r5yXotV/EyznGWPJscqPPx+am4gBwtQQw+Ya9jlY
DqqWmNYO+JbGyLg/0+Tzn4flUTQP19pmn7MndJsR+apDIGUwszRbbGR0KE2tGa3sMI35G8ZIbwSs
mcnIVDadphB4OQMxJdht/M7lHyTsgTR9JYSUZ4KWdhP0afvtKFHj5dryB1jE21XfS5TJsqV6L/hA
kpI4oaczNaB45/euje0z8dkENsl6OVt/+GRAv41uYSCLgrI+oQX1JhjyjPzfipOQ4aREITnlnIbL
sKZXj9sQILR5lEv3Ywi+BBbp91BdXOL1hF3f/3I8tgiiNpLr5hqaKS4Bf2LuKFuZudYy5dnRuSKr
iIROZ0kSyUIGiBZhKaFgYfDeW5lwMGrvKaRQQoqBKLzhNktAH/y7Lx/2KiEkMGZzRtTigri+XyD0
RdiWpWaD7Q8kZw8VuIpHxdXRwpT2a5yxJLPpAVWgGtqQ79fTwAcwl96aPN3xS7km+Edy9pwrMncy
1jG9ol8TUvKeBMo/B+sfXv/3dwT4BILc3e9Fu2uIJ5PWiIqT+fjXpNhGitOctNh25sjBsUI07HO4
MHReoooY0kTyLrruLBFd5p8f8JztV7jiQLmHgG1wzDEk6sYQJz01WMGH8JLFJxctAxLPaIb+9CaW
aEIN3ZMLpQxnMntDOM7sRnCUa4dzHJItOK20v64s+HRrNFsK/V0EiKDACYdwupyCcfN0ee7lzW6b
yAYyNyY/SnuGVOFaZCU0TVx9bmJ3nGKahouSBlV5zSeS8V7HbEXamiAF2j+6YGJa+Oh23NEFFAjj
x+j39+00OKYOQly3uNp5c3laUazgVaAvNPQX2a3dvGvO9/KBStTtN/2ej7Mcw89bQaaVZovfnvRL
42HU5IGtYPvELvw8yuWVX5H73g9PP6/SUJIGBlr1l87IDa9Z/C1faPal1mgUD4OK4rwjDI9vTA6a
160NlM4LkBDArn4covMMNBHy48PEgiSSVOMj9WLt1Bp6h2qfRxcMnwsVT2AJK7xCOp9t3emw4U6p
fqvpYARgwojaw0QkfS9EspeapBp5Lv7wbYibmZar+tqef/6YIJvNNbfFsGE2U3MoUZjVFOuD7Wa3
Ppgzsh1uaI7Ac7pgTYFwmRo4+rq+N/cPsxnfMEqWc1nnq0xslZBA3SumiTIqj10ohWYE9RjYmgVB
Wkh6nr4f0XCzRVJg8OSPiABSDrN6n9IAew0TfEAk3hIM98SWoZ98qm8opwJJ7ulMYmt8Ky2yBoSz
1W8FW7TCo61usgQdQVb6qgcCv9KI5q/OK808xcjy3khi41en9IPhFvOHxusus6t3ew2BrNMxGH6C
Tew28biauNxKavcKfTFYPZmlErBuVecXwlaAhOx+gLRCuNCE2JHuStsUuY82iAnKdW15KGA5fTXG
d9f5aan1vRjT2QzqWAtsTrwHWZ2W4LrHtYu0Fh8XQHaGCOJMImVYQNZjiA+Q7nylx4Sjcsdn9AMz
/AGOcv/80RtIzYHaFgmibVRj7QGzPl3uXvdV80MuAY/G5zhtLryuqL6fvVNrqbYQKaiZeBhTdbwe
gQCyUzVOccC/AcTUW8LnwMEFXe/sYpxc90QygXI2auZtS6JxrbyKg40ecZRw4P2c9H6bi8671K4Z
Tq1ICd2aKhhMdibWRyAWSOZM0A7dK+hq4VmE4EOOVpgBNjXDVkio4tnTFuVZ50H5Hxg6TAqNcO1N
tkk+JpDwQIHPMf9Ytuz4xgAEkrz2OLr55gNIOwhsnLEFbtj48LzX3TyhHSfFEKPOfTSQoPcmKKAs
UE0SqjW8h30R4KzfTHEYkn0nHbzl+OQiel9l5/kvMHjpPAKYpGcMVc3axD5n/HPNw4PDKpr88zvp
YwYXllgqE5S77G4wedy+/SlKMY06j9LFeIMOquBeof9YaYMzG5LQ49qVuVZDNizxwciE7V3b+4uW
rSc/Gft3RqOxPO1AkuNA5jN4JgGS/Fy5BqSJ024qXeyJN+nkQbML5DHMoflnhJT8UXecWZ5F71Av
SlpHYIt+kf6Zf6e6eRBlvu1BvrAvtZx2GGUjMyBQsF94lp0blscxTLKB3l8iweI/ZJkNwwNnzSgs
pKvhZ6rG1xwzIvIbCTznQZa9UROU7/3pbZXtdIX7o16cKk2HxipGfFaB3DiA3R/K6P9gkmEyDMLh
FLkRz59TzFXY/9dvgWUbvRbQQM7U+zEwmI1x77UAaMYw8FsijBJfaXmhquskv2JeSCuWo47uRPLh
y0UfpMekSodvLHXCvVmkjcR828MXABmaxTYs/N+kOLRatqZBugrh9jUsdyTFagXvvQuXGiVcJ/Kl
bIC1YKBgy/M1wLHS7os78W5Yg39teb5T8ofrcjWRcRLWFPk2cXmSpezekXVDG3TKuaPxBKjMcF02
mZXpl7CKeDpsWlR8TbyqivIrohrkwcI2HoxME+k9tyswqpA/SWqgsxyVE2NE4zl7fY3XND04U7Ko
n/R8MyH33KOfRm1m7knp/66bhFI0VAfpLdlTN4sc96m2x7tzRlnp6tKWWB4U65l0/yCgWWs5ZWiQ
n8x8aiwGkd8Ct61GigBY3ybFbiiOBfgsJbjsSXarcRjVBzgKxRWvrEcvJpqbQPv6p36H37NmV+gT
2FdDh0WT6qjJqY+BVJhm40MUkftRIDSG3e5tyPZMXmd7koO3FWQTJerqv4S6/LNhu5MgTlifraM4
LNonyRFnOBpNIxRuhLhHWH5H4gGKIRrO0OqjGZQ1PIEc51GxWFByyl4x5JsEgB3CjLXHNigGpBmy
xUyaVL1BFFo9ssIKbvSFW1srQWQqFUF6J2mF65Ug8drnVDQ6SLe2rBHRzj7tVCgEC+mkUPWfRWHs
q02kR6PeQaheSj6mk4442J1NpivwA1yEEazoZdxXCQHd33SS42Avbj2cJBH9JU3xQbqWQAeNrUKC
m9GYuZ1OH2rqjp/EGF6YzPx1XC8EpUNp2VVsXPcjmELMmS5sCHkeRRYjLCXPaYmKukEauZUnWq1J
aN9rkIRvmspOIrA4zExiP56rGT4mHQ4AnVAkLfS55zai4HNw3kfECcC4y1+8O5RRtpxjUmSVRvhM
bjH7nYVLYX7YtbOtUExt0LvegZKOgs7QX6ICrolWEyYhICBKS4Xg3kR5W7J4zcB1JXMUGviAbxpP
ClHj9ifXH+f39X952Sw7c9iefKV5K9p3hPkP11ZBlUh3u99/1EO2GcWB/UJ1AcsvbUu1zbT/E63L
My9126WhFbSlk09cC3GEuMucl4tImM93k/oTPIMSp6hxtS/DqtXqp+J1mBJzfnLHNaPH8pk3ci/i
cABDIx/SHH9sCo6Rr2OZeK1o+rN0r7EABdYFukWAy74TuhMTC0Fs9NK9Pu92xUsGgeZ2A5c7XtK/
NY7s3E2aS3DyiA2uL8V6hWaAjoJsdL9SAMyi1tHJPZamP5VkTIkog7MFRrlTinPF5pybNMEvVM4h
z9jKr1/OVkgEIkNCWSHi5ViQPucUhxN+99FlqRB2MRtjOKE9mOI/RPKyhP4HfHsVa4V2EcOK2h3b
UZ3y4aGupXPcx9J/01ikv5aSzEF/cJ5SQIzkmt17v/CD9xJfmha4o2JuZIzf9zmjJBwUTyeom++Q
c7Rkg6M5nHSfBJ5fNE/YHkkmky4wRR3sw/0kXDUNEyuX4gessuQQm96ppKiEViG6Rfc+DkGsTbuk
yPCmlkBaSbuxL/1WEpH3qgX9KwxS272I7CEHpOHnWQwebz+4c6oWvZDfw7pqukVok31kcyQ1c7lc
HYln5cimwKvJZoSQytxye0hk4Khi009R3jgZivCLCfwzI0/fOw2VXEg8BqXkPJE6K63PQKUoJs1r
nA2cfxcD2I7o12HPXAn3TJIaWS8AayOnu2iPjFLpKLOzS1VWEW7TDXQTmkTKWED28BLrb64+87hj
Rt0OE39jElIMF9Slof3BBvcz7qKcKXHehPomiHJjs/ULL0YGIZ5f2SUoKKVJ0cwyj0oFnqbu/R/B
4YKG64Re8dy3bBam3swAz3S3tGuAIEspvlso5L4A4FQexa/wbGTvazduvPEEHjAwGamJk9U4lV9F
ZnPC0IQSHYfPUb/0mQMZcOH85lQevIZZCcEsJriRe98Vsw1hBcgSYmXyaPFwVz0R5xm8TtmN6Qhv
WY+ALW0EFKMJoZvMm1D7YJC2ZtdeT5TdJj+YgyWbndidWUH9MEOldBz0eMDiktwpXZ0qxUE/jprZ
932+cBeAi+Eq0Rtk7AYR8Z8IuajQeX5dnEN1WiYZ31RC+R5ALCV98/JAy+kwCkH54wW0TPqmuag8
sS+/ZGfah6P0bQBr6E1/bK9EsvkDr08WAZCOFVWxSq+HbbDGqtdwW2K+ORyExQM3YxQ6BxA+NtNy
6Mn+vL/uxG8gAbs1fU0UaFHA/Y3r67Dy5ZsJGgDBUhBYLVREgRPwcN6p3RhyMMtfkdBSa5haA3me
oaiaawLH5kx7l2EWA1O9K3PM2S7BcW+JOGJtV9W5f57U2A0BL4CnuxS2x/Hm6NRhehf0ET1HeoPV
qtoeEeA5UpFzxzXYn8rPdqLZKCRWNtHKlsVFgUIPxEMHg0cyT9Mpyb6bwwJcVi1DTHLGeg7oI9iX
qD2Zneorj73a0SLf3QluK0js0CpuZ8QL3FtomLgjaupsM6YJNABVKzZZp8Iit3s4qCkdvRJ1aRW6
tycSQJJ1ov69+sH78loahlNMseV6Mqa5hAFW+qQ3ncJF2UEPO/ySoMkzwwE3V9NgIGvcyakBsDTi
+LeqLmkQapnkRXJGFwFdq3mKP9M4YpVjCGtvS610FxSPw4eXpCVIABwwtaBPY41TEolw3t1lp9xW
RSfhVIoAVL0lvRd6m1efAEbpnExCKJ+8Ydd+4O+fXQ5GvoUtpFmo/fuoEymFe3cORtURXacR8Zf7
YEgi8XPNoNuA/1m4ybgpcWXwUWNGwv8APuISba8AWOdyhoccTV9kMkIWjkz9qD6z+AzKljJDYP07
hPxzEu0xG6LRMn1tMwlFZPDj0HeuAFGaxqIWQF46DhAIwOAxKSaHxP4lIcFYqokCOvU2o/+SBfvX
DGd9Tqf87u7xwRyX5HUFv6uLTMaTjv1tqmYu9/7mKSkYXJ/mQ1SAmpFytuYB996E/knvpZUjRY+Z
4xuug2qpiYxlkB++jBWTMuPvztP4IdpELeLGSCdIY6VDe0el+Hlrf/DRAaOZbtVNy7m0yqCD0VTd
yOqtAJh0Gp/ayOiqYWZ3uulWWneDxGnqNATtdBErujob0RctCJLVNEI7JFOmMOwjPWolzddS/b2L
EBBJLpL/7H6BzewFhj7aZ3YziiHATi3CDIce1KsWqMj6KFIoI8TIwttFhMsOyXYKl2GE2nQRutTw
jFqTtZnJNuYCsoqvEXmabrmkrebLiPHdZNTb+TK4Kud2kyNAtgIfHJ1WcuR357VFvDMOqHFXU3+Q
ERzjMDKzVZeuopfa6XJsS0G8unHFSuIuw5fHS/SqcNkRSO9Vb4xIly1UlIN3B0oIqhQyesUPalO3
c8UB3A2TB+Xd4fn9i6FIWnIdmeptDTRT0biDvYwtlm0YvEcJBiKKB85e6N9sA6GjpwnnVCKBKZNC
JMbcavEB4H9Mx4sVR8jzt7C/Y0GTssiCx+0F9E7HMK62HKyIxsIjYXDCaJzVPIxmDawJ4UhCxfqs
ae1t5oxyJbkv6o0RxU8bduQTkCsadF2kik8EeJDsb5XoUU96t9iras3eo5b49qmIC3B57eifBDne
cJMIf2I0qJXWJUgBr0mSBhiLaLuL10ab5SaZrlu6eguy/aMVpV8PFcxcjkkTBS9OWiNf1AVvkLLm
SVEcZ5/mc7TaUAaslKXaW/2pknvvW4bP6qpo0SjwmDbfzOPieEfgprx9HvTzD5rqITZorZhjDvh9
otT4EuPju12TsfTldIWM7X7EtJIJcJEpwb/OsPnXaB4aR5B3yHaP+WaUF1VwbIa2FR8363TLWq1x
upf61b3SqkKPZ3G3CKiCafsOxbAOsJGU7xtWxzlOQHrKb+Xn4v/1t8cX+035dfmAQM/zxl7JDHXJ
S5h4EJsbKlrijHQvbW93NmqR6au48F9ODzIsKE7f46/7mpGaNNYe5uih03T+XSn7FwDSs0LwVrTU
3daD0mK8nmfCz4znt7I+NJxMcbh23/+0UZglLgnpZoBTW2wmWgOAt+tqxDQNfwF0Ldqc/tLTpc1B
IbuS8qono6yzQkhfP1NOhVDzhcS8FPr48fHkfkr2Zdjtxo+QfaA+EPOUwcrTLpTgcgy79wBLXPGt
z0IhTyUGabLj4wwy7J7sf83i1Y15V596WlPNIOw0hGrniHvZZf1qaeK8pVwi4m68ebN9+5kGotcZ
Rt5sYoflXnBai/w7MEnASEtwqfELEjzZrQGMcrQQK8sHqzU99ceiPsv2aDQFhZKOsoiCRkE5o8MG
0GcUs5BwPzlWi9BqQaKYD2gyyspC7F4IQGeikcnu2nUNx/y7EzEuE0WC4g8mvbIFl+v4IE9yXCaT
yBr9fpH8WG31rA6CgnbNlfHayJBH0/m0FnmNgQvLaLDOx8/m2T6zI7WeeeGqXnbbnVeUN4F/4z9o
QbEseaI0Ktb/8j/gl2214Xi8vhXAIgAe9aOIN2npQNe2HEm+HWWNTvTPYIu3qVlFYvsUYDS2TlMF
9M2Jhhph4FzYwOsydW7DowMoecy0EChshkfsh1dme0r5kgntqB2UwelVwSq2FOX22cjiY5Zm5IKY
DsAOqfQFL2+6jqvvymUV0wAI0yD8+SUa0Q8ghXcelxgDneKHaIVfJjJQitwxKbOREVJsgfds1HUb
B0kcdv4lUOAXwFnu733OltDohClgVv8XbU0G7dQmsMdB64AGeFmi2VeYASCwJk8i/+qJ89SDzIl/
E+xDmS73uLXWc+pBWIHYluGYoLk2TdVfW+BQzdTuYb0AsguMNRtcdfUmdHTYlghDxOUckApQ048H
WAeKYPmvLqsDwtB4dib80nlZwEv0CD/HjA7QW/5uP4EBTlXPwSoCx+wopVPitwt+P+lE8DfU8kAU
bEDmH1UclyciwcaxKbn7/QRBf0vW06ZcZaQMmKiJUIsc9rt1OoORSY+OogOFF2P/kGg6PL0BZyZL
cBkdFi3Gm0x/ujbdOpYEDjrCc7kovJOii1zxAPQwzLgkA5xL32jqShQfHOjUcou2EjSFcDSqV+Ho
KG8uD+49pH68ytIfszRPoqmmTEMpczn7dRNSkaW/QYEiJCV+aAFTeguNncc4iDJciEw91NvP03YM
kflyO8bXXuBzrF4/pRO3aXcZ0a5byrfsq7VONvzLkthD/PvnS5RPoP2t8WtYbz/CTwXWxsaWX0bl
4GkKm8tLdBByXOGuKH4ixuP1N7mixmJ9DwWZ8zoNZ3Tk6HMpcTTRKS5vViX2UyL7D799RWWccNG6
968qMgvR5qvh3o024dTH+q7uR/a7Zw7PPeYvzUJbsdnsmvKPAmC/0wV6wIWOLXvTW3DoX7M8EGJb
cvXgmIO6D/jfMUTHsE1+Sh2LBSXKRySgK35fVmE5vxZlWWmxzlhEGckPqdsefyK6dwXK+Whtasgl
z4mliDKNV3zKFhbTO/JRgH2tZAw4Y1sCLk6BysECzLn7QRCg6lO4PMP8xBE8dp0Ma9Y7t0vZOkHI
AnvhzaFiO1OGe3zNIyNxOQrybkp/FDZWZEmxTSZvEXSnQMYaYYRxjgQvU13xYp1QF79LQO7D+pDF
kzNb073LiwPSGYse2M6UZ0RqDQ0qE1QoEnVR0/mJ9e/fNSBcbmzHoP4nfwIx3vLPtUGAPFKCh3ov
wnZXjWOvprZN2Rn1Siy2hPF5mGzuWN3WDgUUzztmr3iu47GRs3XtLTE0ha9BEeahjxtLnycMGWmt
paNx4hnKWubaQ53N6nCmS1zlteOcgr/KYPpm1st2Lk6LC1vh3UHPBPeak0+ygvsmsNwCIR5traoV
LMqLjRbhlthSM/PSR9cqN3t9vs919MutGs3DaSRQZdkEd5j22XxEzV9aemrajHeOUzRSKbxWd/ou
zqu8W2z0xbkXjA8TNHnyK+oIEH97i254NC0RymKZBwo6usN5Qv3i0ZA0TJ8EKMEY7SpS5kTORkL3
avbjbB+sisuwne2pY3aIKumSpQYGeyVJLpS2nQWy79weccIE7c8BGD6As0ozanvVARl5gMMzD7pN
gdVhKWzly/uQokgcVOebaQsPWcklZRZFqjGLQ+JH3qx/p1f9n0Z8Ukm6JhWqYhJS5aHrulYvN2E7
yRZ0Z9s3qDuSokEo/PkC6dxrTZtBZDip1PbXcR8ME0hQkUMTvmxgAomv/TKiXmvDi+f5/tU7soA1
+aTjJRDkfjy/VJjRSUv1aszFb/D+Nknw+S1xylu6XsqmwjEet/BXYyiaqpBXkEkYg6SDJeV0EOv/
JGgDI2hKN004NYJlPcVm5dp6Jq4t5yxexJg5RxKHrucLyRbu5cxg5OgLidrC3iES2HPdvdMVRoFu
3QZvg4eyZe9SuOLmgY96BpVuRdLXS5hx9LjWoWqX5Db45FPapEeVN7nLYC06wee9jD4nGSg7DV+r
/zX+8U2+AVrCbcMftVGigTxJ2n+jEAqOwYtYlBi08IadGRS9Khjgnz2uzQmjsJYeYg7T7oeL0Rpr
cvtFj9xSWSBxY0Q7/1oBH+wknNT8I1CmHBgLi7eZn0X4kV7y8BeJTldw2FMC1kUWmetpOsbpcNIF
Sy5tprsMiVx2ImVv7ROon0V0XvCu/Bl6Sn81s7ENjoAyzpiO0a8+4YLI1vpvc56LlIjbScGK3zV4
fRXi+Pq066zzUGctlaJb44vNWdb/ITCt4vcE10FFyRli/CGLbcxS8VRq79kFgPO9NS2K0FTX1K6e
w6vmrbZRVkxgVRCNOkNqKMbAThxS2tcqjFaUGGhi36oGqfa/s2pTcdyoaa4tAIXn1mrWhIwfZOWb
9WBeHdakBEOnVqzBX7yq9O6lm6h8KhhhZJEGz8zkGDfJwgbrgPSF3K0kbvTYLNweqNVjUXvE029/
WjV8Q4D0M0oECLNC+vB0GY5nMJ43vFY6Ahw+w2c2+6pnKQ39M7l48fCfr3noOmhwWWOBZEO7mw6J
Q3Z4k5g7qPe+VkZpcAzpHOnBsIcCMVg5oZauPiNLCc0QGFxyn35YmRvTkYFm1tsN/hfU4XVLwJ1H
SujhkwSqy2/D32Co7QWQO09tIsJ8nFRXU0GfMlz6wL/h5LLmCI4STQmL1qN1Yg1lzi9kr1jDJ4d4
CJGVrx/GqNWjWVUHwRmRy9oeHqMf+rVJzzAZ1Ytl901WDvlPCSIqsHMeT/13G6s0xk7kyYBxEeaY
47r2mX4gf4cd4tX6ievGE/Knwt+augAfwwHQwmxNd1Hx+5paWut/RCuAfgfUm925RKqU1pvW/b/R
RKnXSfMNSQZB/nEtWnsJEKTAk4J+s/L4oT2yL4Gt/twGb+ZVxc/wNeYcCbvRh3PTAeFet+tQJx7a
qCTiBFFgVx+irQwdcTIredLqd4nUnU1KvOAwEAzb+gPIUecVzvgcb2dTx//5n5jRefqyKR7uz8TS
dcFtd0umOKJo/jOM/3BPwcxNvlWvBDLBVzXjpqjno7JG+2B1tb3F2/84o9Oag4NmrAIOYLp2A0oU
1nNzDpuFbquFWvGCcG8A0DrPF8fJpXx/xFIbHBEc6HBwFHu9gBf0+XWGOoBoOd+1IoXrdY5d6jJI
QCO7q0anPyZqt9cmRA+YGU/w7zXKXMWzdVpiCkHELeyctt76edthFfRWkTaWs4dU4Y1pholkhY+A
F7TcsvWq4eypHLlG746mXzbNhRpYDbJGXo8WSqE+vGMwHuHDbWrA1lZPaqFydinlGiuU++Sv+lQA
ZOIUwfvF9kzpJcrz16gQGe6vQdJSFTSyZcKtJ7YTZafrS/LvvNLYBYD6Gme35fqBgFIIQI+I7s0Z
C5pHycUjpBQoqdPtjNzMUNGAuQYaaeQHsvXvx5OqjOFg01LB555FEbfiMU8Xy6yOMjSdxR7vJolw
FjzOFUkU99ozkzyVpVaZYLwtvtoawkxuvWdYdfQC6zkyQgVFMT/Tknnwc6Rh08JCdw5vo8xSNAnM
/LUmBwh+UwbE2ZACChOdUOql7rPOC9M1BJ8u/8i3n/jJHSNtAbKy4CQqOPNbH96ytUQOTx9nueJZ
Kd/93dGx6fga7gsvOzFRT4zOqYhDQZ559ewmzZYcBF4m1vMd877JwxLDYy6vhuuLnSBNat5jR/Vz
fGdQspnym8bt7ACj+uIOO/zZ37p9Wg8BQme8b68BfVIbpX8Nk2Tc8JPCJ+dBGHtfFm8bbrUKp3KW
8/dOJ6BOSJCnRZCNhn6OR84dITqb9ocxKgTgYwzmChuTgQjwhxkiu6Zl2PMbFMJm2EqEeVwV9+PT
LxvoVU08c/aCNdXFRoLkZwnu8vBUwyCWHOQa+ZEu5mqpWyyqntfRCk+I2YHmf/rdG++F8x0rr7F4
sU7oMIa1d0tSIguPoxiYHm+nfWSszdxENxQZp7OMTdD0QY+LLpLDovACac4+EsGLGlOMmQAMCdiw
68pbmARtV8n+NUFP/hHBRowFE7TbodL74NzsQJkjeoW+y0Qta5ArfqMMTK2vY1VhAaC+DnjXmI8L
MA15tXQsGW+sNythRcCwCE7e+Z2MQovBTreITXLyXa4jeifbqPYqr2IOCbp6IKzcSQu/i4h87oUg
2xwE/E1n/WrCgRPFvlRIi4uGlRndl1NJq8AexR4sMolY2CueG5+/8tUp5bfu1WythZuCOfzaAF64
G6OIOWOj5GJmr/PnXBJZKs8S24pzePKKIlLKu4Mv34RtsOipQlouXtRGvj0KWFZP9UUHYcskmT1A
B0WiDLtRMN7X/dpH9wBNX0r6o9W96vNNpmY3Y+kI7vuih7h1E20h5T6MXuhivmywmL8oaLnEmgao
+ZCV/zp7tu6aISldRBovIiP9cB+nuajuuSiw2Ac3bmrhceTh6eUq9iDoxT4WdJUcn/1pOb2V9jCe
zdPhC+f2hiMWUklNlVwA8/oteaRn3DtUv1Vh73OeVH2ya2wzG9Ruo9aZWIcu+amB/NngXPB4cMC3
oaZFNyiH7Vg9a7a9h9t7o4+s2/PynXP/a7o1tPa6Cv75QrtqgdfJWWKAA4UgISwEs6Qe8sKeCkcq
kyWrmRGN0xK6uakpKM+tth+xJHKGyka9HJlAFU8VoOpvePNCWVksjPHUs+qqKvMP7CT9VcuyEEpw
2O90/2ukqceDj2nbOCgKNAxw8c+TZKfur8NhD82K+uLOXWtYsrAJDYHCldvzSYHCf5QalAlKPA/L
ZX2/xbTI8thiDLiWYsjJqOqpIAL9b5ZiYe4j3MeyswEXWAy4DFB3TyR7Ge47/6njmiI5zk4S8QaF
vO+AShyM2Riv+alnsCS1uwrTCbAfQZZmqmYpmCO78daGa+SdTDm8Mqos8rGf5H0km/X7jZ7MU4Fz
Xb8cR+ng9BdvgMVBlfB1eTA9FUbm9nMUiYV5ZjG5m7t+iw/LUnqIq1+XLMXHjkoU9iNO7hLxmyKT
r/bJ7b9L5otPf/hJqLMOiegI5wDRveoco89WtQZaSlruz2VTP3FwOqm3yBkabiDcUlYMhcClAGji
9x4YwVzHP8HYr9p3VHu98dR3cYyo9cuBp3j8KwgapChqPcC5x0TMHM0U9WBVaZoW08DZpHiXyOp3
IZ1uBf5gUsl/5kWYxlcaijB4ZkPdmn93TKvC2nHfIGo4pvJ1WJcrtF86+ydvZYKdsQGA6skblRki
j0h2ltqXYaCjdcVyvI7FBZJTbmZ+wvBT1KOn8k14loY8VjeGW02PvpNF4d+cJ//QBWQ7+caiiqOP
mW8QwtHrOhBnLnapjWk23jnVHTETBW/mgKqbq0uecEY+NBISXBTkQ2KMkbfSNyxbLYUzsmh+qSl3
lcJNwJlo50e88mfaEYY0DG4dmprJJcs9nvHOyIKWLJrDuoW1U7PDfxyHq6kkVTqSKji89J3dC0xI
vbv+SqwfeSIpQdwKXUjVFe1Xcvd/M1cW4kwBHauqlBxCarxzOb4VGw62GPmanvQK8gksEQG7ONgM
zcGjRd5gqt1QwCFHcTL+Cqw7X/Q7kUyUg5KDObSMAqTGNlVuYj1OCd2OmJeqB2miUthYFHOqC6Za
17auMmwMqHc7DJjhEHE1m1/aocjBd8uKr1HMSiVt1lgmI0MnvKmFHjaTXmplTn+UZ1zAaze+L43S
CwFqrucQ7bk7Dyb6RHW1lKvMsyI8B8HdBQ3/GSozVnZQNGkTOcXuXTE58Nt943g7dJfzGxEHo/cQ
4YMC8apfJFnCGvzsPYxtE1qdKSy3EubSiKYpBoz6z4zT4sElO9jkttQrnfPbnmg5wgVXlJYd4fWe
CqgmdATCx5/X1Mtf9nmoA3DtPgIPPFi1IBVmttU72gNvj/9lJVp5sgyBaJfe3U1VUO7bmOAhy7/Z
jM7Mm6wS3PDmS5LSRJ1CXcYkslDbbp8xh4jY8lUncNBqDusNWWFofq95Uc9R+TvgB8Yqf5no0Lfs
88vh13hc3UZUsSZlxVgKTiQzi2ei3Kuv56e90sH4ObVldLBaFBJsJNLkhfr2h75rhJ3hUHHJJqDj
W+lA1YzX2csmBnQXWPC1wDFcuzdu9EWk/HJDoe2UWEhm6djVSxeKwAKYuY/6FpAfRbXUIG/hBchV
rTPNkAUPzkkdXjXrxA0PSCSgPUsz6BtROElMD180zCDm6y+E4S2B34huSiHFA9PQIgysull9bwVY
AQ7P8wA2TT9VJoR05G7M+zpvDOCmeOtUa3BselkzkSbYf3C0xUheixefo1kg1mjdFq5jw2d1vAbC
HX7HdiN2E+ZIzr6DeSs9MP8X5ASXDAZ3/xU8k3aFsH3HRCNiIza1siTEZvTQPIGxRhDvbM43SlTF
Cqidd20itKz1vtSxvt/zqampPbUBkcxdaObEYZjDJdvs2slef8dnX6hFzX+i3dTLd19+a8kuFiP3
xXatr5lMOc+lNnQ3JeLUvyiMpLGYK75TdZHZkL0eUgETMtUp2iJdyGRe2oIHA/k0LhqBMTZ6xC65
SEBVjkdd5URykwh4qGR4zOlW+9qQEuSY4jUSybyHbXZyHMW6eP/FiD3A8W5SZatT4j80jYhz7w+g
kA4xF6B5Jq3Ed6ufuCxx1uLXxLnWpliXn4AG4JenrGdpbbKIc4EYsmD9CYxtRP15wfMcYJUqrptZ
jyoQzOo1vff3XcWDdkSPwwtRKf17Rdh3t0JxUChKLib4n9m3JfqlavvIspPMbf4LmMKYg20r3Eqk
nf9hU6ygvZWk/OI+a6CrBQCYRyI6qcUGxxUhR1NI9zCWfdUoL2Hr8ZvmIRDmGUoeNvZnrzQ3LBR0
P8PzAF3jIo+9nKHyDgaQ+eMQnv3WdRz135ueR3NITGjc02Of64/R4vyiSEEoX907EjUBvIwi7oKq
SXwBXstgcqrGui0HShCaCvRrdF2JzHqOxUzx7UTRVvXzeGoJQXb3Ynr10oXyE86gN3Dh3Y4HXhTf
8HZa3xn05yU+zvtcvhBmLG8IZ5FX2FNt0O2bHVM2uj9J6yvhi8qFL1WZlrqAQDehCeyj8HcAT8uG
LAgVfChfloO8GtHBZ9+A6Tjjxms+5d5vMkOyqD9o5kvEn1vvjuSb0n9q65u0YUyXHtk8VgVzvXP7
FsHXavqEXdTp1pe4Jiv8ggPpr19G/iCwJdCZw+K9kL64YcZl2wkH8vm5AygWE+yxomPbIe5sSxqs
ygPWRCXHHOhbgvgTST4c6jhJKtltCbDctlmMgKGHMX//w24jqEneKqrVRgu3j2Z2LnWZOIvjEySh
lOru9JNy8KxYmWfI8JhFfE8A/ykD37W+qC0TFfp1ud4kly1T+pJFzAgvUM4q8c78ODXBA4l5myj4
pspIZUkHtg+Of+S7Joi2TuQywLa/uO76PDbyAg6HSAubCpkx4Lnsy1QRhF1AiDK5ILxlqsTUQz4v
qbC49Pw1+be8/mJnLwly+nxfjqWeHrjTeS2Xgd2tVBZhdrLOkJD7zK96LbBPSE5oLmLrjovCFlIK
OaC+bGygPdmAyenI7pDtycA8EAg6YYtMLSBQtZJ9/YSNTizWNMlLUkQhDUd+X6Y0mSUFqgxuHuOW
MiCwI5JTxfsYsHr/AMg+C0tkVzoynKVQF4eO9+0T/OpdOrhH0m1m81ngPIUN0tLFGnQI5pC3JpCV
geAD8h10cWe59AbR8idE6PMTL3M7jIEaj/dgx2yIEVyqeBrYeBVvPizIA1CYR+ImW9M6WtczySrz
yHTbtTTFJVqjnash3agjGq9b5zhV1CxDtrmNfQLuLcmdguN+hIKaS/A2JbzTcscOINZPC9vYU2n+
YlSHlYvjYr+XWqV+78kRuCyVPed6lxrgkhoXwM7h84UIHEk//5qU03q0ka+wq0Xl+YkU3mBJjv0E
Vn70xeqOJ+r0r0FPVs0W+eU7z8G6CHBLEI/emWr8gknDQ5QBriUM3fxwBp3yf2fEbQC+7zzvOcDe
4wuSwFWuomFTQF7zZBwDD+Eb52+/8/UvvBBVQb7DXhNnfGb2ZbIcISFoIPb6ogezq/0xoDZqdtRM
2hEgq8i84GLDv7ReaPURlvmy0CapZpzOpCobOK/XiIm8af8kEDnkg3LvGpXxIfUa7rHh2B7J7eR6
tMQmabaXXGjxaoCZGAH3uN0lta/dEmXNX1UvhbF3e7e65AM4XPS3Kw5ka9KLP1uucl1Qy0YdfIhH
9zxYxTRTeLYvMfb2r9xVytuW2L0INN+OSBcfXXzm8krCVM4BSUV63RP2SL4GXF1ZyKlIMn5KR0RK
1XwvqJa3bQISbFwomY3ek1yPvCvJTDjCHOkNzz+/LTtV6I3oa09OQ0J31vLE0HeSzIeTS5snS/8a
9SOOcYsoGIe64RXS1a7yl//DIxJMzTqgEqunsYONSQDtdknIzQHEwTi5Ml5x+hp4FGYkJ3eyWqPH
PAyBiFPUjUUAOc+Xe3WO7IWfivGgShT/OqgUHAQ4JxDy2ONGA5uJ8s6SJrT8+BruDSUVTDtUid3b
fP97hDlYnkZH+vx+/3Z3NXqUaNrUGn8Zp9uFpxw8aT67tuV0aJoWT5kWhrr6ecFZqF8XmbsQ/Rdb
rVhGOepEaVuWgKA46ScbZan7EHOzX6YmSgW2XF9K2LnX7/3fc3Jo1luEtBtvLNPY4KjXFkfVqVOQ
YlaaA/40Y8B0mJt+Y1URNA3kf44/I9Z812Rq/3nrLbn12BRghdzZLhI0ywIoOzYkcEhzhey/ANDl
a2YKU/GaN7BDavyuBRGpr7wlH/zZ9uMpPYDYQr4icq2MCUj5gFSb0drvOL9dq82DeUHStMc0MCuD
TYrHM/szlv2EBfDhAWajYC9L6MYVawXw0Hvod1430Eb9lcPbBDuhLf/eaFJmrHsQif3RVZYqzhJI
u6qe22Ibvx7SwWRNPD+CSA9ZhAC6gnnlDW+cRb6Y8tQfA5RCStfyaLW5hPKq6TOcKC2MZ2aezYrF
sGantV0xmN+dDmEFg+/8HvLYv/JFmjKY5GDoc0QARVPZ9UTngPFHUsv5FsAuTCfO3aGR/d/qBTkd
V72mLDkMIAz09m8zDHZ1kd9iGR+7BPh6KQpcLo7qzDbhnind3vcQfbygBM3/0/WVtw3jDUSxEffX
Yigxnf1WHRDuui5mxlxNiqncpBIFyJ9mX7+fhz4yBIo7twDz8XhiHSMpT3nVC+141VVAuktWYRT+
OK5kMP/6kJiz7/xOdcKpjKpOEH/ZhcKcr75oCT598n5W8PgsUgtAGBeSSUStmawQgZQoPx5kJZ1E
cZTQjvZRvAhlQFO6+w0U3Ev/rJ9kSG2T6veV6nDPRxP+CIpLmYNHxz7JlnJYQ3kdsTYdzH7oxyAr
KsEa+MwTez/pI4Oy2nlALfmoH7Bo/bWC+v0qAsrrkN49ygBM+8lgbLBLzhY3nhiu2S3QKCyDWaNU
RoK2rIktHLOfrj46ZNUVubjCoMYhX1y1pE2UVPllbqfIfsVXw81NdkizvFTHZ5CgKS5UH84er6Eq
0P9cKaHfVp9/BZsRwqPgsiNHBmvcq86yP+pyhvubUTTSu5Qs0VIYJtzc4GqkWnYaMluR7n5R9Zpj
jNZukiqjaOsotkbPsChNorCasTPDCyroydunIMXWPjqB/JRHjVSsDr1gRrJHHDlLRA1Tds3llJTL
SFaSzwrUvJgEWHTudjMvdVURJ602ZqWABk9geMLURqKDpc637UxQt0/aZG6lcMVDZqwEWy34r7O+
kP+38orqoTaxBCBWSsmZUU296JS94fMw02SZdcw387acTsU8nqUtCaQLxpBTDEvnxkHLZjG8ND4Z
efpp7zEBbvndvXO+QeijiS3SH64Wk1vm3BaxkJEcd9odjsVZv4dcQkG1sslRcwTv9OCX1KMo8EaU
1/BYygCDItkWGJIz86oh+o8Efscig1F+55TctGJ2CVSeV6kJ9varCZtra5u2L2AqIrNHJC4gNl8M
4rB5lK9YGPp+OpGdcZogCsgqrd/1wJIAJ1C0PwhtGuM6Z1hOUIIOaccYcSd9O3xF+eM63p1PoGVX
D3g3WUj6S0xt3KeJxK4XNH3oE3eO6MA7xZB1BbFtvlSRlhwHk6NH0SU1nxbRN1UJ1Mrypxq6yDWT
ii0Up5xp+YyLRmaB0geDU1wwtJ0CU/pQI2m6NtupgBcaVuxU+vketk9++s6U1ZHN3KZyOniNhfQc
dAxgAc2B81cQbDSmUmteXULcb+BmBcO1+Zyi3qTLYbldmVBV7aEhB7aU83ZruIdJNnDE/Id7YQgR
v2BSDIW3SHPYfA3asR8rXUTdLyEVIIpaiB/o4p3Bvwpttg7WhyUimnMeQmmpfoZqGkYtx1Gz4pGs
WzBMvIe0OroyuSql6Iqnbp2X8y2+yzOhOhIhbtlvp87MTYr+dkNtSCOTy2qoldrzZJGdk+UnD9jn
VYjcfOBsr7/irTXWrDp7qVUbHerY3DAdjam1UCTqkvKf+WFvvC4Qzhd4N26uUZjnOW5R7J1ZNDKy
XkA/693M6DPO+Ht8EZUsG0qVLtMhHq3BLxK8L9KPlHG8elbr1heZG+bZwf1L/DfbC36QpDPyxaDI
kCda3iGhlVQyjrlCfChbNqxkmXw9LXg5q0AUP9U0Dkk8aRGNOrd2bdpd5rmu8Ow264ld9R9ppFb1
dPP1hweroTNInCOc9ubQGMrQvhlISPnYuJpK+GbiUN++briedfXECX3GyF7m7kGZ+sSCqWykA12R
8L1aWAFBmjTogV43eO3Cvr0yhtvOqm/4MjabMImlD+xMT0+3qDDUrELceK8MqMaDhd1myUbdCwFT
7QRvj35XxogNClGYfKoYZAzgWCkdjGvR8zR6rJfCAZE2+/kMBw2lh6CxKrf7CD+P4FKsfFyyoc/F
SISBMZIPepdEYPQ9ZlVBlX9lxebVDWlXtaVBqPHVFjh3uSYHraNuGD8VS7UEO/31lxfuaNIGNt5z
Ic/UAyQ0p5HmEvvW7/4cixXn0TH2NpgSrH9I+v806cPj1LQIkeKDziIKFkhlrwwN7lOBtp3vO57F
/X/ildHNatMk381LBpS77ZUktI8xBuHYmBZuN8vmUxpf466d6lKCddes4JT/hKgg46cCENQVT3JE
XuCAg6v/O9AeEW53QYvdESNDK/6ZgxMU/0x0ztjtMcYVLHzHDmWW++el1hTSD5Omy7y1hi0rFqNW
IaplNuXJT6hCDdUZJh7zKxry1LOPvPRxOUsKKnbViM+5jDwcvvC2PvI25nMl29Hvb2KnodinSwHp
D+ssKZwjslJilAx1funfrPviDLfIGttsz965JNP+eBAhDdRQvgmRzGuLndtlUwMk/unj1f93Bz6h
aRmi4+wQF0YTzRJVJmIdcJGXqBPVKj4VjBkXrXv3r4eGKm0h5tROV3p3KnJGj2fnnvB8t11CwIe6
rpB7V/jMt/L748nNad9n6sR/o0GGQ8LC9hvWR0tpvvBbppVd/zvmaeYqWblNY2cBuczRmaeUhG11
s2g6UwAjeHFjSvNMfvzjy5bSn0YLYyyrn7ADpBuxx6RJ/1m9QIeu77/Dp/u0EifN8xq5FXAz49aj
GyfhM5veHs175WgamnNs9edK5QSAbYG6zqPZXihNvhm0dS2udOe+Bs1Hwb52iwRjvJ2O1TWSg2DY
fUaBU96cng4A8akcmuY8/QDj99+84xawVoLzZFZJv1NK1UqLT15EZjkY1L8W04zpfgnv2PbsYJGo
WGuQDyIt9/l+YQYSkyeQyYuBqvMipllP/h3/XeXicBQauaIC8TC+tCW1Xt813MUxB591HH4mWSej
ttVMQwW6V+ioCUjt4YWHZkFc+FsV0xLUVhwCpfDEhGALB1+E2hVBGJAuIDxshTECjDe73bzP4oVM
o5woHhqTpCqMo+mJFde7NcxUxfKp3ZDwByE7HgrdvDlETjwV7PiOICc9I8JZMmTNCZHpL51Mm77Y
QEnf+7YYil5XJV9UtMQJE1mE3bc1KbpPnDaDtdz7+6CTi32nx/HLysx/VZY6cJZ3vziGWTW7viJ7
sVKzwFFcFyPdah4LmftopW47gdn9Xu/ZAeLCTRl6PyU/I0AFWKucnjoHEjz5k3yjrHb1muC2CheC
FXwuI8UVuOqLUuC8ikAyJlMFP9C56HeSMHJuazao5xzKxhfFhzqHC52DJOv7KFGgHzzTVVJlz7Et
SdSSz0eFyQz2AimKbDRHONYgizYdr3HCm1SkEreI2cA0joEBnOUp5KAJ1oJr5rMm6JGPRy08Fzvk
80C58bVjO2UOmOh7G26FiskjSx2uBuhAHnw95xm1fvVhLGZVtUpNUuT/LqVjNo3o+LRfnct8pwtj
1xyeYh4AKwitProOcnHqqMvkYpFLvy8Cm0yPfXXBS4d11r4srM8XnnNEcGkW4jRVFcc0cZ9eggud
wYOIh2rSO6dEzwNmJHwz37PrYMGoyy8JnUCHvRnCFcXyBZdZQv3JgEFsSQ1JBZE0lvzB36czmCiI
s1kBL4VHgKW9LmLAO5FGfH+oMe13/O4f8jnB7Rdd87uGNu0S4qrFT5t7+EVv3Qk2kzrb/AY1Abw5
SYUJASZfW1+OkNp3Hzwi2C7oBPE9/Y+v0GAYzAaoXXqJwFQ0rh0EdE7wOouzmobnb4BLJxsQx0Zg
OxLtqF/WvUZNj1Pe5jFJ25AUoYaZJEwQWf1WuY11tg8Dv4namJo/H8GMvzoLFqo5EBdYl3TC9n0j
0ZkIg0JY861OHF4McnKP/j9gCJtHB+kxcCxt7Ft8x0mMamAzoi64mPBP1ZLybNUKsxu0Reg+jlju
QmPewupq/KA4UQDGxeJqlfMw5cV5nWapQm5MTvcgK1OZ3MQt+rrr1xol2XlJQVfs79l7Pokms4FX
GWpuA6RgngkkYuysgcIRCGn3eHm1oG2LvsUf+zlRY+TGGlbyTYkhC0RZxEZH3XB9cN1qPO1eXy2e
aoB8awXrFxWruUI74XQd6079hAFZe8pCUYmgy1g3o02J7pFBSI7MCRFIEk9DcaO2f4hPdwkAGsnp
uEqJLb6u4t9GldEmXy3SifPZp7SayF0Io9+XVW5t7/VD/L3AyUoSZvmWCGpkHruge8Xo/k/6pTVq
saHM3E2SAuTBuPie6OJIsoPUo+Jh9nXHYsorL9BQmcZVLmT0SZUCYQHJLr8qCD6NOAvEHilK7FQb
y4qOsJMGuM4cohqvca2ZjoQmVcFLV/hpt381Y3592Vh2k+rRBOfPo7kpkxwaEXlYHk/nro/XgJgh
7eMi8NLHKE6rkCZSSmMdriEfC0XaE25Rx+PGgpU4SgoCSk4Cj2FjsZPG37lCelOIJXql2LfXziWk
vFQ/2TG7WG+5Nrg1Kfv623tb1OVRJ3bj+cHEeerBZvlbDh/bbHm5EncaTiwJx98UeeQR2vfwo9ZI
BD6sCVpR8Ft0Zyj1rtEOs+E9E3mMIBsRMY47r3wAei4/vdVRMmVNNwvzeOAUZLM2CwIJWbT0OB/M
IFtEhFQ5R1IjSRh4lWBwk1gOhYzGHejQ032XrSWNpv6l+PES25qDQGiSKElKosm7PLeoQj62Hkit
9vM9ysjAr0C7ljHWfFjREzmYCjDYZMEsSefmpwT9MlStN32wdBPrta7S+fya3C9DotEYbFy6ufAX
s9dzUHg2fJa6Ef1Ab2uvIj5ju0exBN2IjpZvVNA0Iq89eqXs3B2vCCSpSx6E4WOgENU9gp3kHnZE
D10rswp+KbaozIwar75D0jL+ukrjZ1njuw+lCEYwhVXiT1YVaed0PhA8ebXD4HKcVeJH/X/oHTOm
/dw/efDrTFAHQF4k+eh/E/yE0ZQ/YjyArwny+HW0AjTT0RKy8ERvD2sPfxQxevdMMgCGJZ8eFL7u
3ilaL73tfCqs7/BaAoSyVPR6T6d6Let2OGmNHEYrPnFmUu13hqbc0gP6LYqRVNnA9+HtnUDmX43R
v085c9eIQTVgZou06k8tLd8PbQaWkErYFIlCA00FiWxf4CsTYW+errYVqp/vvNRLpne2PClCB4ae
bj8qUs7nbQAaAgvRWbFznNq1JYqwhylWfxETK0yT5NL5D3dIinyOpeYX1Wi2kfk8A2Rl/5lPet+V
FI8gUWN/2sxIIy/wGbIOB0FsIlvrNXm3N3/TioELxm3mn11mkLNNc0r3pn96Ow3tH6PERBXOKfsC
a9UgraOJWQYN3ij9E9tRZVSzFKknUah11+MXt2r7K53HpyqRwF/gpzgVLPHUCDZYHzq6xmX2kSdm
vtymMjEDyTiWNF25Mz7MpQm3k6QklrtCP6+F0UF3vqJc/mJGwwM4vLzbsIPeM7TottU4rQeXwTFF
XIwaQhkno4tNeCeG5jphEliK79yZjYhFJNdeVk5a2VVEAJzHh3tLKjSIdC+riui5pQzzDdJZjuPK
sbmnqw56ibVOfMgh5BeI0QbEKni304v3H4r2CiKFXo89tJkiwvIKuV17ka+pc0hruo/VFs2ukD+k
2U9DLagq2gUB6vu+sv7jQm9DUyZlqzmlcbKabo+KTNJZsdyf8ar0sQRUXmECH5ReLFzQmaYDNNN/
CqEw9M1gdzDoJdy1MIHWiWP+BOwAdFYLtYsDTbX7Y7zVlDeKZzv0hN3m5KQ33sZkkam4Hx0vWtcT
m9QokAUiJnSsTrWnRkBNjWFztrwA4G8FHOmIoEFX6jqFjsQLKnfwrcwutCGgwGKWxOZ17Rko/qWy
dqm0AJ494KvKf2U4WG8c2c3nj9Fm5StlwNwZuaqgbvOe3oGBfDDXllnIbUc1WuP505p0doSr5eyw
xf9lDtnRiRuxsYlAyNzWu42KAjHZZ44uFH80kwcxtROntOsGcNpTh0b+4Bfb+x+LfmAbxMvhs0Ig
LUkNN90o3NnulNq10Kane1mWd5VA5M9QQQcaKNusMy445EvUBvhWMNP3g6aRB7PNWxqNmhcegZZ+
YKvJjxecDx5pH98AMe0jUVrRxzKHb8ItrBWi5QVSAXSaM9cf/PgV5nS2+qL9jBDlmTRuR7+2bsZT
i8roQXImbRtz83Rg9nH+LBhVaAC9glEAge3XxpMKAnRLxOw0qIGxlW+xkt1/RFTnx//XoQ+Y+sEP
x0f4nS3AJ2CMfV5ED/lB2h/7YgtzMMeFZFfaLBdu/FN143kM4war5Xtu4LQ6TDFqCehy/0wZKZ4T
plR6n90/INHK0XtXbnW1EPGEAlAVKfmtiCQpvdYBW6cNskHC3I6BNi4aaGU+lp/w3WSuAvWJnqvS
tslvMP2ZTig7aCLfh3jZHnH4A4G0UqEzEv0216NGokjqq5f0mLo7l+UyUCLYaCWcFsCatFaw0JpA
2vmO3URok5ylyxnu6j59JVKTp8XGkKPr5+ycrPG0487wvt9FXVQBLMqlIuMk34Oksa+1JDGQ94cX
OYcGUnJSuAsh+aiXvOkPPcVu2uZKztAy/Ms9nYOfstndPpC21kCc3IKegihrQo7HF+alqVQkOQhD
+w52u46Uu8VSYhNa/dGAeGfZNnvzdJ6iL0igSlVBCza9gFF4cMOJRT23TPiGKGbZcC6yUoMRym7o
EeQ1Mb3G5QHi5Dyf2LZ7uUoiUeHGNfKnLmebxxoZ9sM3uUiG9uA07W1u7Zq9Vwdj61LiGe38HLV7
aAEHWlw7wTS+YBk7Yi2xqFGea+aCE695M8LRD3yimA4OOoR4wR8QwGHOjp/64MTyjyI6ir0TJNem
YgGTJqSKVFgl/3vUKAlxfqGbEutscOA/hd6Im+5Mm9z98ZE6M3SYuIumAzcysfKnWoVjJXGgn4/J
YgVB0vnpUxtHegene+18tIQgQTdU+E9jXor2HrAFm/8/PE6amU3dvNoRq7tPQ+A5ekHBZ32qXCmV
5Eui8xX2JM9fMEH0mRt5W4UK/r+8tRvmOO1H4KP9iVHDRNqNjWy6stdFYIVF47Ffl1dFRtU7mwb7
/Y/zC0o7jf3/vngbQ2RwdGuRVpkt8j0eCc5UA/0NfBNAPEKmaiPfNNgEbxM3CwJ6zkogOZ+tYwjH
PJZNEXf2u+LA4IV1J0rr9NCQzZFeUYDg3W0wlUtZGmoqDZmlisVno2iuPt6z8Tv1J0RWE43LSZSQ
4Ke0HKcBbVlIPIdfBqEoSCdGjhYIIddHSwmJD6RCwfkEP6KVczpZUw/GoZuSJesmeReRhWHiM+Yh
CxMU/jfaqknbkS0rAwSVDzid+MoJRveLDaceNEklwGz36dEqlB0BV3NwquXuJLKNGL5rcfi7o+wF
HuO/JYCkJY2zj4PIURiG95LI8k0deKX5y52Xwb3J4wHqcxS4XB79l395vFMpdg5aqZ99ieJiXdAo
o8tF9Su3AG4ZzzYhKzl3tA2TdNmV+fqxHmwXCL47T6pUTTv6o65ubzF6m8Mz350v6mrN8QjeLjZ5
y5M0ZyO6g1PtoTBDbaacAamPHxho9/4qNcPDlj79OriCARtP1G2PQV2DbsTAxP3Iru9OlYAD9rYo
39MyKaD0ZNR5Wxn1fbIXOYHnTAgApJ/nm48nPPjUXv6lq/YWH0je2Sl2bKyV8o7iSWsqdvhB0ME1
z9Ay4+3lmvgH0sSdeBQAfiMHWt6PGSk7cOHNMWX1vldw7gvNNjNADa2jYGsyxs17lsgZi+5v1g5L
tXdIiS6kQSS9AluInV1hKdWEF5fPn9nb4V3s+Folo1C3iuGTx+43bR216rvnb4mwngSzPBut5nBT
Iv5zBGx2bapkIfGNp4yVC50h1aXsUJX4mFXnQPf8NUfCYihaIe30AiYm0R9kW//VN+jvE43lGY6q
cSdwvcTp25JUBN8yEh3f8ZzqXfRvSNQaETVlIC2yoOXrS79QxnMxEqRav2qoRh7V6QwzNbwk0Jt0
nJWBXWa0YrLpDLXUKkN7R6GRSZw50yJ3jJdDm42uojtXl8xPvCuYqtcLtuPr6aXUhHnQD/Ia9qcQ
y4JSYfK2/tKG8/rUM8Gc8UvZPknXZPLUmE7RHI+55RbXlAw+aak55yPLVzbukpf60exEbvRpfu8d
SSw8sUf9bwV9r2KRZBp+y625QQ7NjhRckWovFB4NiGxA2x3/Mn/DXxv23BOStkkcleeMQq6pOz7h
fhda9Z5k5qP0RpL+vu2AaPZYPKbe+BoaHq1eSR+AGPJMqkM5PwrjxFPXXijQcOpdLIpD3HQaRa1o
P41O6X5hn4iqf+Y6MnhFZ3j0o2v3ZBRr/wMG3b1kcH0tLtD5jgWPii/GkefWSR1Ul1zd99lCjd9G
OKvLdSLo10W2bS7+vHcoNH4jET4terDvzHdMAPXOdyg7OnuwyofwFn/MeN5yHjV4yNg0SVtc+EUf
YIQJOELoiI6ER/zZgV9xQ6cM0cF5g+YVwfBXLjd3eWpjHOA2uEtcy6eGtmdFbWC/gX2R5NqDNzCf
aZK/PiWOgXx1KZFLprEA2VLkUrKHZnN+jQDd3mVOyVLCvN6gcCLWofXuAg2pWPP4Hwk8BRylT9GY
wHsVOhbJ458ULKA6rOH68Qhxr0dbU+qzJHiudTOmrP7uirK9O5sPiGha+n6ftULvcn8Y5cyHivtU
dU9t7pP6M5YhEm+gr/vCLglMGdW3fLnJmfInU9lwWXPexMXlccE+F7PjNNMjhmgGAgYOd9o/AKib
552RVVvgQWW+EHIqeBL4D2STY8yvTLQRz8wBdBR60zfTZb+9laREQw3aJVfOill+l9yaZ+fhqruQ
EanVTLaWKpXeDAjb1nLGiNOcBPoXB/6G4gz1VHFtd3R5aHu4i+FS12YvP9iBW08kvAXJpBOoYV05
W9oij0rNaAM6UcNAkEYhes0m4nyRIs3CcpnhmgB3NOh/1FLihRwWLJ4XYUWSINLDpmXT9zS4WeP5
0/jkEYpP5sUur3ZUyTardbtLIh8cwIESvGCp7hG/bi4CbNLnRAHAn78JtxyvFYGBAhnrdPvI75Eo
MaPaU6Gu4X52Dz0jm1e3MMIvXxVuTji4+nHB3+aFXTr5RiQTsSjf8n5wycPvqQG3DEPNpRrnHuBg
BHDQyNbA2l6YiaWkJvux/YIbflNvFRsqPYxUWtMdG1GDG+auBuq9Iaqpr0wGn42eDTPNkEL92RHI
kcxzR3KefQVRoqA9rvG/o318bYGITldAftG/fOQApLvLWeKmRc/BrFjAUcspOj/jbBNo12wtW0r5
2Qx0dQAAaWKEqZBYT2QQe9B051ewUezYTPK1w3ZdK2VfRhCPHopK3L1P2jTDUdW+LMTdEb9+MshP
sFW+WWgN8+3NH51HUGZ6MPYzauPa5OoFK9obSg1dxdoWr+gBV1YeuNzxFZCFd2k3sQihA93wkBR2
u9tl+BJMAqqK5UoKJZkEYC6Nbsj0/reE6V2w8Ae3t1Ov+xhL/sxyB7D/pbE4NwYIGNCM8B8lymGK
MBPU1hxAA/tIe2cInR3qw8xanf7HXQ2ZIRXVLECPVAjcPQvptVB5Uf70JaattfgElT/k3YbwXXWR
03VeSeAQ/+MosV7+FXAKcJAaUyaJAVf5tpfZkzTu8qgVYE3RVI13QFWwa3XjF63HIvXfXKcz8K+Z
J5ihipwzTiS79HqvVFAfpB6nfXhgzmIGcuuAhr3fjKoHVXTFmtNPnpcQk60F7N9t5bMzk8vvsr1H
/bO4/IxjaNdv9MX/iBJqo0WcbKQwWfHM8GQW4aRrPlh1Ee056391LcQDfzyZgbdsfmTOiqMpSIiZ
smzjCkqNPzak9Y4nIeH/go94a4+C7sO3hC/zlDQOxH4aDveofyczoLNXlCppqQ6zFlb9RcUggyj0
8Gk/T8Ib6/j4SdW3bptRDFFrZWsvtvXQIA7RYvoOEcqDwqyaEPtA5bQ6sPfvGvXqiJz07ecLuZdp
HdoqBYZAihSuZicGBTh2TmC64P52W31X5U8Zk2Frq8Nd2iGsFOdCi+RcbbXpnV0d+4/954hWfjYL
KaDwPrQzAd/Keh+DfDD+cA2HcVqhu07Wu8ei6AP+m0d2gDmVhxw24QhCEDy7hephpriCXlV4rH3Q
2CTl74FtRRyKG/tu2uuwxDqDla/xG9fNhIL+NQyOXOdTUrBC3De3ucHAYT71+2G4Afj88vcFd04c
wjXOX2Yv2jAjHb3fymnGjGWqZAPTb/X9pQ0dYbZKmJGuhXllGrm1za+NLY3ijab9zc17HFkAmCQJ
HX9v6cE/oGWcVrDStFpwoGv1qrp/kk741rJ0l/fxOd/Sdj59ybBUSHpi/rRr0aO4exmY4j1+AnfF
yfresWunJPevhaIW+8+GgYqntJZkgLKjK1pzmr399z5x6U6XtQJwx+ke3fj8vSvLFELxZ2q8CZiE
HtyNozJ586h7iqnDsmwZ4mioZ+fAp7Fs9sKYs3QhwSH7Vh1q+M4YH4qCkU+ffO71PFqMcp0J8CfC
o2vg37/KD9u/SZimzoH04DKeldXf8e8i40BFAVMGrnplOMGF6i3FyD0Zj072Dl+d6//9DcaSX02o
zreDNbh9N5oZUpXjmpyaP8x5mV1bhSm+//zHwx1xqlM9ZLhydD/QZZRrDd6+mV6bAovHyqn0QmOL
N05OqkOapeAZXoTiH00X4ubhNxhsYrs+FmIC+BGlCux4l63Ym3od8oG7flrXM8utvrAFPJaH7CAf
zVdu23jxUsOy7y1pl4nH0chpAzNEstDCsQzLe6vzboZEyG79+WUdr8ljcmIolTfRAzUxWIRlgmId
5o0ySZsAJSWO720DrlGnQPMa+sjG0MCjZot2ivz7hQD1OCQcLuEmTenKYODoqzAutMVqtRwI39m9
R/K26bv2gDslkna1TPvFEJXJTbm+ntcXi3OZrfU/1gbjPOH+BUblybo/7M5Jnf7S6aUaWQm9JLWN
BmPDKggI19N1R7UqIGtI7M1SrC1+D8iwKBSYPnzVNyPoT5lkDMKWc4aWZgCC7YjFGrxeRRESEMQD
NzORQxaiLLxnB5IiNf7EQlC1dzeUBTdikZZfJF2a/xPTgtZy9jUhxQRxryTxMT693t2mP10+YVgo
vvYuN+Z9/OfiWwjuotRx2phbyweTUzitjeJ7ck1pye7AvvD/pncFLxZjmnNjVPVqhs+y5+A60wMS
eRQByrT/hK6ZyFQT3LxN/2H3SsLirVXUbPmuuQcwfrLgYlH39yU5hloMDMoS1CyfmqUg7hBx1u3w
ytEiJv5L/c02YzEiIbQPsb6QBC8ehOxd5gjBsWJEJDxDZA7MCU87Jq/PpdLspzU5KecDmw+SjfbA
e8018G20+GnRWyx+AShBezfsmYt7bTDJOxh7J7hvReodqRtxv17r3OZOChIrSJMhSPR15Ten+0Ck
CuSFmMdy5Yk4JUzAcsRMYTSnLKZlq+370fy1cgD6WfF5xwockGIFL+XK53W/Lmzvfzzr+cO17ssk
ieu7iZIyLCI/3ORDiwvBcZmOcDE4ZS0Zs8MLISe6HlrFBCE2EMP8/PP+/RrxlQoCZWsv1eQKIDI9
g0HfNW6frdTQ9OiufWAgLGMB0pn5OdVV1Ydvjz0C0Uuj7aU5pCUAmmZKARp7t581RQtz06qxT5Lk
tEuh+1ogAH6e1M+lVluJ3Hz08iczARQuYKqgUvotDl1jTNpoHYkPqHEjqJZgTy4GMjUNUk8GT1wr
CD8khJow4dyRgEdeqH21N3gM4VfQNvNJelG2QEvDdhqJJaZ/Z5O0QXpXaPsL6no1MZZcok/U1GF+
vYfNxglCFtcKMdUm/kDSVVveZM4TnHpU/mMl6X/K/K8gpt/KIQIg35gZhB5+wNsObNBxvI/n9mWK
7gQ7I2G2z4AvFxlReqxfDmzPMGgEjAoEPNPRxAlmhT6iRB1+ZhyFQ4booSy7I8pcChUw1AdVYYVn
rjjFwflhHXGPxGIUhZ5FYT372CQfQuK7K8H8cbDJ+I9bMKO51rcYKmm4jIyLrsFWLF+f/GsdULW+
yj8bO7xdWwG6/xJ3ip5YkV4lb5dsWT3BW7cPaOrui4PSQOPzXVmVFNEsMOOBHM/fEfzpm2Q6DpJj
wILhSZz7xRK/ZL+VDiWQ0Uldc8iPkoggpaiLOZ4mLz1FQy2IiiZSr4qlyiAMmuKbWA1NcaFgFW5c
1M4bJ/6nqJLo2YN++++kUqNshXF+QrbskRW4daslDSMaEs9KhCdByYSRscE0FiOb0H21edgx/LKv
e14M4Fa1UHodOYdvw5YO9eBC7701GxAtoq9P5onYCudf1LkZ25jVpiZ+0njrYVK8yBL0nweIu7l2
jkLqkYsAUV3j1d4z823t3vik4nhXh89fMf6Miwyt82F9MpegdHa6XVH9aeEVMrbty+ufBtCofCbd
3dXLRPq0exHhKyhCEVYXPjHVRgSQQlhHzjCauNp08Q5k0KTigIVgwn4OFjROome0ri81ixsBfrzR
KsGMYG3IAb+udS7QgpYkefG+m6EIshQ+2N5iyEBgItRCul58gO3nkXzBd5KwpClc1A/bihaA0VwT
F9MePM0mA5jGHbON/npYQFEWzUk/a+5ruvZEQgIXTewkbvnxVg78OgYSEV9Pgf8WOvXW1AFZrhbn
Bnmhe7w4+hURlZ/EukLsC5Bg5oBA2DruE8mNsg2wxWPoMglpAWhxLGJg5ExJ5S0qK+qJtx26v79F
Cyh6SaW2ig32GgSo+0R5t4yfqNeFGOY5Okf2Rl2JWRAOmfkn8UwyAZbnetCVauDP4lT6tZ+f75wq
jFckd1YevxIBZK70pAjE8rtzmT/sWA1/BqoeKfy7VtV9IOKjbjMXchSml3b9TKi5nSDcLsed3fy7
1Y0cbcpWdwWAAxkpfS8njLFfkG2cRDydxli/esoOFs2NzG5M2evlbVbuzGudPbjSvN4IBVWd4vHU
HREnPyorbVj6GBK49SurOmmS5a9dhfoyuJ3taCdGCPIrUmkZ4DsvfTr/N9fm4MufcV9+wuVrtBYf
WZx68J2NSVesy5uBAK8SvishRklpDhfElzYfH5yUgfJtcPR7jdKuFLDLtXLgrvpzyqmBTtDrTKUL
Dp79uzVHSfa3CGed0R86rxjpkaNlwBMfp77Qcmdj0zuZ8o7LSSvarAs5QdW1bU6wozXQOWjjKXjy
HSdpdiuBCwzVcxdpWqvyOd50c+g37YG8/KXRYfMZ4Wunf7oq4vmcAYVfvlObl98oDwcLG9VwLtG1
wmI2Rjaz3E9178+PBR+ButNAlbHkOCqXFtmMCX1uthkwdcP8Dw7fs2GFI/aXVldA2wuA+z8sqRQh
7pC03a8VjJn6wiQe1k5yG7WROqiF6NVZkgSsR5E6CijwJbUmZ+/1yGDBMw4GJrsB+LDZiGKYEKeI
mBsVll4qhuwkV5VEcsaqfuAtSHzREiuqYo8Lfi2CmB0svHEhXLgD4y1wJ6LhMn6u42ozICKS/2Yo
7a0j2Qf+4J30WRT+SBgK7AvNaM2YfxmIbdUGtAkMu+fZEKfQJBQmlr9QFF2B+W3mJ4bDVTM07WhY
HmXmGAePaFh+2vCtGtz3BFsNbB5BfEjFpxUFt0uq0hxXoaIMh1FJYLwmGPNdIxqnsteDy79Ae1X5
/8KTHGLCoCts8zsuYsfeo8f+s0mIykEjBD6Zro5vbrbAIB22rM5QvFhItNW6sxr/ac+4WrxiV4XV
1TkY7mL7yvtR25oB2uO5juZ/pgEwAMBPjgs8cq8vHLuWzpVl3koHb/pqJaJ9F8GVH/+vsHJn+LKG
m1rqzLnhqZQTJLOYtFvE8QNtUk4fdIzz54rDr7hQC7xxcanSqZTzK9/RUf37ZR22VY+FD0eBdPeT
BLBY+DB/i/6yLqqGmeJoE9TwTFMlxQKzP1qeWaLg06NkhCRfzVxG3pMafyApr0/uMrkW+M5neI65
1b3GB1LMNeTFAAVDWEw+fmYLVFZEltLXJoQmrRIBWwrOlX8iMrR1UOmr/8uE3CQII0ZjTzaQNUbe
wuh3Ff2UAi468ugd2aohjhjyAT+VG76YOkqoGwWdYfsFVQDT//BfQCAXADtfM86VUh7DUdLP1JrE
Zcl1vXqHrNwpGCMkqKsJ+DPztkVeEQkxJPvjipgD/l6SUaFaXzQH/NHkBFy2icF/ApgDtluBQW9P
T6bBp39kqjRarsy6ChEvRnP2U9FhjRYWq0EPJE/KQ9yP7mWDbF8UA3zpo4kMUxYi6zHgunMfmysN
a5nB2mQmo47J89P9ydkz6fKRXXDqPzYh35MeMdCwmJNWf37XLnxJr1D5ZpZ0EkkdQ6U1Wem+FUxi
jAnKAmmgfId2YN6YpR8jmDTdCKjUnoJwmDe8oIzcBpaIlAgFpC+0YzBwscMEJMDsr80wrNP/rub9
Py0z5D3lmQSjqrKupnQgprxR37CBVdCFCGUjoVBlA6qmQmzMSpOGxvFqc8x0stQOC5XDezPbTcf4
FI55kNYWI1U51Q8miWOGCpK+wQUr0hGFfhbOKl1PItEG89ow+kk7EP7Kq2CGx4gDFuc/rZnt9vGL
uekbJspNgKwJwTEhnh1vVRldPO3Am7zio20KfEEoIl3tyY9bJJ7w2473GsPiq9FC0RyH8PBXYtZe
eI46YwOzL0Lv115xtqYQM2+gwwsi5prvGa4RT87NvmApxSRRowG9B45yESemLuQop8ZWTrAVyYqg
lF7xif2Um6eb4Lm6lw5u8nHC/cyqr7zsqZNV2zEK/inYHz2+rqFTbMWNgWLQQUWiujArklAq5dqk
+6w/3qlB51MUMWPNStTf84sOI3uXjCWfan1kppwnsiPBrYBpxUZb2CZA4uL/T9eVgWWgaxlpXwNb
huS7lb533h9pyW9PxS7JrDFqRRoIFihQPQ8As5LFXW6ISmBcJAOi0WJy4t6lWjpeVzD19J/ZvJUC
duAfg99Z4ficlVWc2Dq5qBMITCgfnV27I+CegwRpVPD9uYxVu19L6p4IjvR4rvJ/KgZAKGKr9q/t
KDkNouLo6+Jx+V5KftJdyt4VrhmofxqUDJVO5YMPth8lEuTP3tsG2ZkvYnCGGChwYELtS3PfXjtd
3FPJJ+s6Rg7XVwyM1VsQm6JVUKBx1wqk+cNDqy5p9Tr3F53IPHLK1IDwbyG8cvsv7ll+Bn1CCIJP
2adqrJFNiwfoYQczfpRGteozZpcLNZUfwC9hr170Lk4WZjNq9Cmloqq4hXdKz+fTioBc8vSSUJ2Z
rfrcdjZp1QTFBrUFOS8bwIsnorf9BmNEEwtD8cvmMJqdadAWvbx0F6cwUTN6zKCu5nUGdEgrOWp/
10CnaVfIp8hFWGl3/iClJy5kHhtVxsRTPxDqzYCD/C5PFD87IMF4PQTxMPFBQrYeLDMvWws0YlXj
/Y7TY0fwz+naBVRw6Gxf4THKP94ULV+JQNe8HgtyISX+CfLWljVlEIazC+LmHRvTo6zqfU+Z/1y0
HsTUQUtI3di8+Rp694YMBAlLktGAljd/DIU9lsxYUHBnmXr2a4TUJ13S1JG5+bkOUIuEAnxPK6+9
9IcCwQTr8+dzUVyc2c8Y+MLSLM9D5YHl0c9vRaMTuJ24a8LsgPrfpK3LUcKftSlzV8xRKzFRdrL0
XxhHajdqlFFUPO7bTaBSnOy3d1Vxeg6jDGRra+utJM3CJMaXlBlMXoQIIe6ZXqk3l7cBKQxfgj5L
756JhugVc1i9q2Av9zSSzXC1efLks8//dKLwQevLD8b2UhzoJNFZ+8xQNu5YzntMiQDP269u7kDE
6ybSfopH1ARagp6+mIb6uDmo0hVrED3SxZspz5X44TOA/x7dLGvjHVEcijROjQ37dC6jtmw/6wmY
FprPVVdaACZhqM9p90v0LMRqql9B+QC7pxDo25yCBQ4p8b0JityfIiehT5XahOwTrNxCVEx3osex
tI36NkLNBE26TcSHE97hOdALlxP31/mPsL/kpG1Sdvg+wNhme5S8fsoiajk9k3CYyQux+kiQFxNG
o6c3jsqNANyWuWYEZ3cKX74kMvf0VczLSqGyhMVpl675gSiq8xOkjLom8xB+j9y69d5XE3o+Wg16
klgXM6lf8VQkcBRWdkzcGVj/Qrh+uCABRvicDgOCavFqLbnCt/2Y8e13Qh6NRv7NDtc+mBZx2t1l
v9mcWejY116CTLFQkALibRZPabVrefCxog39P3+uwWCOlV84s3aBKljscNmS82EyskE2/sUurusJ
BE2Xqg2kmifaPqdKAZYCmAKdUJJdX+sESMoTtUfVGkJh5kkKSjcMLJGHnijDPZ05uRsBYBnFjkgv
sJbFwfI2tOWZoGTRGLx7RHpKnO4mj+egzhdRkQBTppJQIfCxrchwjkPfdhEczgQ3Q0+gWeFgs5Pj
O+92qceGSm1V+3Jv9Hd4luFj9KitaQERRfnvUaF6ouWU9/bF24L16l4KbohrXEOUMWk/IE5dji6S
Gi4DnqIlRUKnPhzUoe4wsc/jt6rmIDW92Edygj+SO87Ab1kjxit1d4t6iIqK5PSibWG9IhRjVSG/
F69/Kts3vA1SYNQev1d8dJdsNVHbFApgjRd3ql9wKS406Rk8n/hUnpVIVGxNoPk8TnnMzsnBoDXj
pufm/6wHDGYsChHL4V43EKlzL3+aAxbSKH11XPsfsCjT3+/5HDp/x1oyPgDhvI5/gXVncWODBHQC
Er3ZRwEa0ogmCX+aU4cMmkBDE0xf9I2EOGPxq7Fc9+c+tl0SoV4XG64BAtnKAx0JEoKjnXrBjuhB
n0zZoEJ1wMlG72hAJoY1ifal/IPGh2D/kPYqnTXctz34VwvbCjGYHbkUWHO5axNqKM3oBPzbG+1r
jz+MDQAiOWZymVW6obAs798Zl/a2Cbf/AnjocvwuRLHGoc2hgMvIZ9n0A8otj24pkzmtt5xaAXzR
OhXFZUjAgn/4vbf7mz4XdgkyoINSRQIAJBv4PxbLrZbLQyBhvmphkcfm0KVS4sCO683BPM6qPG/f
OPK2ZvaBGjW+3VEiA7Wj4Ng+CErCX5BR42vJCyoO8J8OIyAhftIccfrgx0VJH0FsEfzA/A5pZS29
1Lx1aEtICRNjbt3OoO0xOKileTPZXipUgVBGWS5gqhkMCRmKzubzoiMjrXpG3GD6VkWM6r9o2NFD
dsagKLc+GNe9izIRyrlwkjJy/wVbHzK307NEteBzH5o6Yj59Ho3YcI1kvvlL4hJFznCva2NrgTd4
5JYuN66IOe5KUSMZ873LUf5BaAo/Th0s0BlW0FH7F8r2tV3mS2nG4RLlZyD+9OB95YKcdt6aBi1i
+ZPgmzMUA4ZfknRnufbfldaN6dSmtI0xFLpz7h/qZze4cnWuM/TkBBuTA0um9jkMQyUB01BhWAZF
UY120mRQt9UAKY+0EVbWlKSGwl9+wl1G1gXyACdIXX6krECRxzzs8QVdPdW4Qna77V9U5g1cCrJn
KN4480epembwg8rAjVNbtGaPXeW7EgUB0sFdfCLRfaYDx1b7+ERUuqaKwKyGNJURCevfHgRsUpkJ
gicIi29/EkbnzCa0wQ0SdfSL0KeBiTF4qgK+oYXugCw8Rrf+JEjpcN3olJG6FHBNlrPRi1atBlgT
BbXhTwKapVopraf2u2lG34N7hjsD6PI4bADd3DnKbZjSeKf0ARTjZBtcnYTjhVVx6PnnAkTqZKjp
WxKvWOBjaMwIRpFtHwRzJztr+hNuNHnDAEXdceMOkXBUOutNFcbms5Pmnbzh89zxiJYSEGBi7LDO
n0tYJsoyRQZs3knAZJ1QNRQl7xbtO179ODxb60gE0Jh/dAmID/Dc/468lo8uOLayNMyLbuUZozwT
WP3Z7vc6E3pkXb52l6yzlIuRGKmX4vVFB79Mt8RBSw7i0ScPMY+TY1FZubjuNzyKChypFx2f/jlH
HHpz1b+JXmxYC6SuxLfFBKM8hn4JTlEU+WWa7q206WX0H+nSRJJ1bE+1/ZqxiKkJv0pQ6ftUestZ
V7sKRnxuRkxvfKeSrHral9XxiOuTf7UQtAi8t/8nhe3nAwgiV97krOKg7aTc4CPJdHGeK8ylR+oE
4G5z0P7nwONQz+lA6KmTTmqMX+ggjSBIArru+ZlbPg8ANwyl3MnWiSLgcM2fMyUrsKshDPHHZ7FB
WSxjs3pGUPa3TaDox2Bj6f5kN4SjYZge1GJIK0WrL8p3SQP4DP3iFjCeekg82W7XZI+EfbjS9Sj5
6INlxgtikGmMX3G1EScooCEX1WuUgsQza6f8MKgbzKKjfQUUmQ1ib5LzPxSBpijUsjgxW1S6J/p+
PFK/0OcKvXe3RqBODYHS43cZxLe6C4F/ML1AIdInCTJ9SqyUOtplEWrtWOfwN/EUha0R6c+45z/Z
IM4zrFBomUnVEIu1wz41W3dRxt2YNID/ifx8QKn7nRBYzS104xjzAzlX6Uh+1W+snWkgG2NgRdus
5puVVMVxIuXsQVGd420ASclUSD+blmG8rbVgnVEz5ojSWN8cgpoU1jZehRxDZ+rnkaQHnXYm4bVt
3gLzkfz1wo+6K9dJ7UsSYeE2Ko96oI2dCGDZ5sxFOjgQEEdHrUsfxTVS5/C/yb6Jf5bLcHPYSNsu
ccSeB/ukuq4s2uI7pA08DymNldbm+o97ngeahc1tErlGrrD/gLPVv05rHcrxyUDsuKxAAtTHn5bd
GwZq9LG3NHVxIQ5bRTr3sXsadzA4W59Al2sox6Em6Ueu/HUPJxGtFlRL9o3Tk+cb1A3Xh6CsBJPJ
/RAHBKyH+kzNGdq5suDHU6PC8S/RO0PRcu0OqmTpIhKVSpRU2+ElVbwIVXHsI6nTPrCF9CjV9mZ6
fhLsihB8mm3+/vDpo+4fk5qcAHHBOvLUokxzWtDdJHWDrH5xOUIF5D8RDJh/AjuWDwLYxWIcO90P
/fjabM9FsKHINnljUQbe45mqV6BOAua3lCVtbbTz/VVJXtTG8Tit/E1ZzDoph4FV4kdRdNePJjAE
82Sk4p/Ro0fKBzlEjxHAMPkzWgKAoigQJvMfcQbbbjXMQLe2iN6bQKsvpj1mfxUMeGriHz06EoQp
ZLWh/qn60pZWNNWYLefMsgKMQUWz9o++W75rmrh8Lgj+xh0C4+pFUNgTFdEcp255Eio0dr3z36tC
AA9HNmfeNl/G0BZBWWXVhtsL9EEzCjBIrvkRsa5uGlrNi6WhOxIwMCsG9Smt1nvU8jUT+T1CVYr0
99aQZ/LNNOtsZxNbZ/7j2UWYhYW5HC16ljqNCRcRhALUtcke2T8/96eWQNrlTQtIHqwvKqgYxs8N
FY9TuclONPm70PwPNhBUQN9WcwSuoD7qz3hvwmSYimQMr0C9+kpHNyha8Hdx0HITHKcHn56Hi4xi
DFiJ7R9XbKObBez6cN15wsm5SV4qURjLBVfY1MKDUDTHRb7osuEqlRIuwc2Ur0Wypxe4d8Quoi5L
SYE5V/vBqZKx5/UyA6MIm6DVHAjtFNq0NubyuOGVMmsTFXgxZjUTFq8OLWlbD+oDZy8TjT6U68O6
YWBgTmjgamcDF0fegNCWA4Zzzy1l3U5EkcVtHMYXdauWJO/rWlyDrsdRQ8MPtyq8/RErqUeVlQdO
TA8AxLbKTvsiqrWRZsVyXgj9qmT5O1c9d96dkuhRNFQvb5K1AjnT/i0XIDHewvAo1vzaleWxowvA
ASMCZpmqKm8WEe28uJCgZfaqKDSAfNtjuc8Jxq5XzFwuCZ88b+Z/nMt5sk5PIMnxSn0gT/H7GV6h
J1kdhd/9voXs6NFd8fWmMbzeIzq3SZ1eL8tNOEr2ZocSvgsffhXYsJi5u1W3NRMDazIhl9dyArN5
6sGl+7nHg7TUdFQBnerKBQ1ZzcLo4vK8dNqcKMDdz2pZaQakmMT7m2r0Vnt9yrnw0GCkCI/9IrUA
gjD4EkkyaVGwXgR57ETc3LR/gjXDzNeW0vUjF3husxiKO+2o//Lp+ynMcXSTk8bucjD8WNCskYo9
OsRUcsRxU17EdiueHq+oNw8N6lWRD3QUSgwvtCHl4K5C3aOaTz0yYA58jOBzLwrg7gQK/1fVv5wy
yOMuTbcVv66/qaqUcUjmBmHEAOwwXGO8ZWBoE72fMAcnUW7BTbh7YVDnNzyNAzNBHxA71ZDk0RYh
ORDUK+B+TgfeABSkSL2pkO6o+QqADrlo3rxYHOHu+EwY50XpwV8Hg77y9tF5zXFMOTH8w/WPZ7fS
SMkAC5XnirJdh6FMW5MAuWsHIoPmQeBtRp9Wh93Qk6xWUbT/g6qMXy4KgOT85TFXRp6vFlS0b38L
s3MmEIwfSa+WWZq20T5sQvFGNYSin9jX/uEznv4jxKKlgAOp97uCsdUxkS8IRRLkxqXMwGbIzuJR
QOzcR6rH0rPlEsl913mnU6EZPmk2CyexJwtsddjCNX+8Qczkq3NEQ0YkcDnCtnYAb6vFdCpXphY/
OjuvjzM2++FhSAePJVUiJXh4gOvNyb5ODN3Nzwcvf93fkQiMHRBubS+GsJzcjno91YL0Wp4RGzcf
gq3P/pcXBJDKhivjhjXhlZ/Vu7/EvFmkyG5NnJ6cYGHSzTF1YjEAfCv7hcEv4VGPnWOp/59Y8HlI
8HFci9gWvY0f9N4gBKtPvu9WQ3LLAwQvJOM7N1d30nVoc62v4VHvfdj2e1GoxPX3ntdwdqbBc/Oh
xIWyZg8WOO0mhVPbV7vzBs/AtlgqJ5dqHq64dIJyegetaya0fkv1nZfiL92fOvus9HlCZrAE5ytG
oqZPBuomkJMIOyciYEXjYDJF0Jb4lqWdnoXnuhozZ6fqugrmsZzaGeLWfmJ3FpiTJrRC/191SENV
ewPIH+ZJDu8wHZRDq8u/pJ5XhijPyY6G7xUrjgveNb2C6Rkog5f4B5WGcjim+afB4QrssKorJtt1
sgYq+BtzZVp/BiXYTtJkYFj/wpXtXnp5yGk2+wq4MbheSbzb0pvvcpYVrY8pOtOzQJjM/MCbVAH8
t3/d+lIUK6Uu/HDIMkPI7JheCUHx3A2I5F+UfTt33CnioDkyd35LSRqf+s1RpqRhH+nwlYCiSGHQ
fG+qcB3lD9KubFjlJdF/NUsZY/s3ZCLmjzIJOYKh7MJAHu1EPSuMb8oM57oLeMHWiDf9nujWxTkN
Rwf9jFPoesnhciU8TeemD2A71a4LBBbr4enw1889XDqwteBBMyOwaEA5irAdqg1O+dDcTlICAnAk
jm2oLBe7RXN5zIIIFDPrQt0uNvheVtvHTRvazlVib1DKSspyGj7u11tmzqgZR7fiRPz25MTH8NaW
T8eFJWY6A+pXe/2x1cl4HmgC1T1l6WM5fnyvT0Nk3gRwjk/Hx/HFoxmsIsR6ukSDg5cmbTg5QCnH
5qMzHhkrWWw11Gx7TOEUietL+dKj8RvoZ1DiTk0KcK5VWCv2pAkB5x/z4wA/10xuxCXb4rm1MxpA
SrSK6MfoiKheOFF7HavOIEl1DhjPFQ7MVi49JbzdftZqxzmBpgCOgsyqT2c3bMGPBqBuQVb2/aQ2
jNccq6oYAEOHarDiOfFF9f1aSFLmuRFokcvOpHCHfTEaBsp2eym1jteGfyMCnEvFM49h52TUaYYc
gYYDVgu8W6atozIZMSz3m09dvi3l8TPJ6fUVGI0Pv0J29R6N0SnvLYeAh7XPPlLm+JlIDDhDg0uY
D6i5xA4tdI+F9hoDyYvJxCxabBPW376ZNlb363th3OPJKllr0FKzaWh3xqa1NzJxkAVoVv/18A33
WJEczPTHE0M4b8YTiMwo6foNRwdUDIzXfQmBYtpDE9B0x2gcxjD+EIz6f+ojtcsWwm52RAW0GaI2
H7u3AmW7YjCqe3KwH560JoDwjJNBRJqpIqEU04IZjntJL7HfDPjkZQqbd5w7FlOKTsu6cY7ysODe
2D/5vDjIcJWh/pYd9Br80AmaIvnIn7b96KChfwPFGR82kFnE0FB3HVLJgpKj1Q9cKD38BtHpF0C6
egR9IdOx4ec0MmjUrDdKfjU51r0vXJfMgObfQSWe4TVEuBiYrFTBSi8NX5/1wE6oI/oFpQIDzTkR
Wwmcg7/kNVYIH3+7zXQrMqNcLnote5WxYZ5p3+5Ai7/Ope2AwFLuz+Op978iMfGsVMyH2z1qXf2h
haKySEq4GWYUPLSS7AzhMcfTbIaK/f5Ts4dM4bukuz1PyG2zSYz8qOBwrGZgpMGCHr1UuWoIxQuV
EtsZpd67Sz+qS2b4pMfYTxg4a+F46+uFAEJDyiUoqnLmhRWNzBq3yTbtKI4eG8QBkbDWmNOT5RW6
C5X6ikx3y/4y/+7+PDzv8UQoSYt+lc0uSmL9jSXsIQCyb4WYsM6bHxE/PCy3JqBgX07cmvKwCgGX
JItbmxcklhfjlyUvNR8UWF9qMsrTJEG+hctPDBibr8tp1a00b3Sx7BQcqkMbBc2AGQh71NvGjvm6
hVZtmgNYYPecVk+DSLHEpulwA+wx3AKu33s7YEBCE8pfusAmTcAvTCziwr6cEB1r5lN/hh5mU5K/
ojlrLDJG3vbtHaNo/8gdrj0N8KhVgXlK1t2zvH2KlKYECDPg4D+0MSXgdSXHZrrQrCGHQr503Jyi
5WO2f++53VtYrKRWOU0BQor3YRt+fqkfe4OXkQwMY+9xz3+n4QSLhcAbjGIAAi+lyPc5HHUM38D8
0cBsUWk+ETDqx6HTrhmujwAu/B+aVIRN+gdepfQPS7WvZlRLSa8WWdkuF77f8N3XYsNHag9ChV2O
Wcr0/ZdHdxHU50LTnd+3R2CQ5N4pakCBPCYL7K0EwNECa9YWhwDJWDoZdVi6wEqMaIcWB20mefp1
PhgS9p8VqKngo6sterS4mH/eI42LjTUVpNQxuIjH6fYMHZzyyLrgnK2pWm+tzttwvr5i0YslQFpj
v1KIAe+d2cm+qFixxZDuei8DrdUZYtaiKZSL4r8f+nAZo7Up2kh3HUNLU+f4E1B21AWMazMdStSp
pnzFSFDXXMnqpAMmlu/gFk2XM+q1sByUmYb/Onm3zqYlIQJbzPlCj0+vHu7BQBV241VVzYvj6tDy
/qp0uXoujYpdEX/yTtY0tEddSdC8+2RnRMLIR/PMv410gZiSh4YgdVWJCET6HbQk01ySmazC3y0W
3fr3joF2ghwO8lUat/Ylv8hrRber2GfIfNT1OesPKuFxEuHhWr8oo6Lo22ivVjE8QzH/YHkG5MC9
lJNIqbLF5kvibKgQLA1GvySyNwiBR47ULDXeL9bWkF/YVTLJixmDk74pbzx/tfOS4wOOlXoyHwVo
Xk13Tbtsw+oRCL6ARJ1v2skgLfPisYVuGaZJnsEO55RAnPFt9ySCymsqpH647lxUCNlfzioNL3/B
ptbQrJytHm1ZI6eV9jhZiHyjeapLy19uBqaUFncIHAwIGpw8nUX0rUEN8iprbeJzQLRZ1ELp1cIS
QpmusNGi9Db90Zr1c5aeyg+9nFl2wpXj+retP/Onuc+3Uu+PdIIX0nbEDDO7PVZ25IPezrICxScy
ntBbh9ZhGqq/Dq/E0+kkr6hs44XYnWv51A+883IoTYyjdUipQ4d3txob+m2/bEsdDRQIBo1vthnl
xOfZYEVASPCIa6yJPdIp5sKujsV2oo6cOuHlQ4y9r+E+olSD1uFvyfKNhI/jpLauPgAqoSkJ2tPo
DXShGlN6I9L8VJIway0E0CipeaxChickXQqfB+oGoKkiuJPBSzPAVJQTEcoIMA7Bk55/DssO4Thv
rj1bIElkAMdxorlkoLvIb9/v7JqLi8OP16kgB7pr5968dXPxuWDA8nYele/CKnC5CeeFK0eDrbph
GuEpEYo015Ca6xrQr+a6zQGg62htMwvCaPkE6hQIuEqvakJ926vDBgqjxPkUnetAf1Ja2d76oKwG
a2M/Si7osFB0dMAflbBU3p1KVbiRnA/O6a4vKtu2ijk4KQmZFiMsYZ2o/BPLl60dsoymogoNmojU
GwHy1aGOVebZhgdSvUFwIKGg5AP92xA/2Dag+YCnHWZkBVnLnXlM6k8B7M6JIGWdS4giPgdZ+iKs
R6lxWEg0c1dipc0PtO6iaBWru+fbYdDA/Fa0wHrgTlYnQEv64iM5KqxHtUZNRexMErSHZyYfS7Pl
W/cXGicjvmJHsLMarb8penY830ubCafO1tDlofFhdQAO2QG7bVLKwsUG5XkIsvMYtFulcSxCohjm
3qtew6+60c+qAlu/nVxOFeOQDlPY+8fmIP4kjPtwk3hr/SEMVa3xsW14gZVRp3Tb83fE0UtaFtvz
AZQCAYITydhoyhjLtTuDL6VBukYVlrisjiNGng2E93cru9aU/NgsJR+lIJbyCSS50eoQrWOtjbZg
pG3rnyhvIz2u51R4EaY7O6SkKOInffE66Hr0BHyw+Mv+xUBC5wwWP0mWBJYtxXRlBwY+mki8snQG
mwCa6UHnFh0YAarSKAVYUMPP98SkL26ABdDXUC/CZcz3ajHLVFYOrVZ7li0Q4bm8BngqfZBo4TFm
JP9C0I2bXTs2Syac6e2nKYCHxmTqVHUxOHAqFXOQ2eI9bv4LlvZE6Gd4GKrcLFMlooRIDNJKLyMx
OfzAwXdutr0V9NqTdhcBb7J4YM0Dpe1B99xBUfk4apveg9O8n1ZKmzAiprC4yeOovmbapi4/vv04
SRwUR6fLWSj6tnTW4SEOW1SWSqndhQXdprH8PtonFcrDRzlHPdJDXi1HmQ2pypXbUWq1zyYV3h23
IMSyprARzQGAbtIC3ioZyVxK1Z+DLOwNHVDUm/yFYAn40OWSvMJbzHOJyvPRjsW8zp5LaoXB3x17
HbFH8PibOIqZi3wgXa/gNAlM3f0R+d3HqJjhzopdhadbhHF9YBX6yNYlgnlUjGf4y7WoDOS0UJmW
x7iLFoGCqE9zaRYWSxWaSiLehs916SXLozP7S5hHtNibWkUinWQeGIqtuMyAmfMfgJLEhkjESwUr
c3eFBx4rxwMTwcERTopv14lLDfo82ct52d3Pdgu23V6cnKiFxaRCSEU8EfSvJSNy/ictlOOZYw39
kgXpiMTVrV0d1q+zdUd3vMCqWfZYHxdM/SFFq9of6mrv3uB0Wj9KbT9DPcByF2s7Kld8XebJ63Ho
EcDlt8RfwOvt/KYEMAAtWK9gOH4WO4vu5jR0eNaoN9gLgZdSkzVmn4k2SBO12xknMhvVUssLwcXg
vNsQBDvzsciZo8XCe+bK4YVoDYOyALTDPL/cT9VH5pgFSwro+WoVOf38AXd2S1RiPbTChWfb2SN1
pXYPiUwDjHo9BtCNiWov3cYzqAYl3k4/Kb+H2QkO/q+/IhcPCz7hLsGK501gFrvLGy6y5gots7ZN
0fexHger5fJwA21khAl9FhXgjnB2unfJ5ftK1C5wwq2e81dLggbFJMAMD7jWHO2AcqdLDq0vUlG+
2n7wARJ6ZgWQoh06S+g/BTJPGZ+O6XVyMuQImM0/KLb/6GgaLw2JKyW3CGtq+A4fWedCz3CUe+ew
unt8hpAVVNIhAhM3Fv9rmCPnyVlG5ng514ONEoCwMIiTtKf5JCTJpZaklL/6v7+IAgpou7CuAy9U
lM1hNND7T7Urkb5csVi+fhWkCLwPgaNA9ocUfw/PUqJWNGO1dWiWpileDPdFejnp6wh7WIxtinU8
grRGRmRpI2cHCgSW1VkmiPjekRKYxQYFXetNNsVsPGi4jFryaCaYyQqTn0FDS3SOEppXd/gJ+V84
vfhI1h97e95BMBs+zhA+pKdHUZUWsD091HwoRS96PJ3r9RbcMA0pYW2VYTyOzLUer2GHfN6tjjCE
rQZTyCFxBlN2eiBhh3CSQdlg3/4btddyBehGPXiygHGKOCp0llJUcnwC8ksF3X+48fgRxIdKmN9Q
71rK/fT9I04dSEsT+qPN98/Y+Odijw0L22pH3IeSBNcC4fLtSKvUyuj+OzFMkWCMzRwJBuJDBMgE
82ctOAoF5mGPdWshMGsHT0j0JanAJZqd5/RRjadByTKd9MVV+0mJC/ZfKAg04KZB3wBdkjxzS4vB
k4itIzYmbASWrLSI2228F9Ik1XgD33goSZtVjzsT8Qf/TYongTlO0nVtGGiI7J2Lsyo4i8FaYOf+
NwKXUdXw98E/JZZTZ+eLfTMAQM2DqZekuMdbBzK8ESqIijR0rj0bR9rV2kXk1iYawf2sPT4abjtB
VcWn4JRx+xKWqSCPLe32lJSAvrGPSVQaXgc20zbVAzAsZAqXdOR8qdkF1gfxtXNlMZ0oQt9Z2r/5
MewVIhTzffOm1QiMuU338173nplTlpx0yAFLYLbu6hTyJ2cMPLvRfbxkjKPH6qAf45QDmhcUU5Mk
gctaEWFiu2l/G6/PVYh9MwjEch9XypFj3lbU5J8kCI8EslNCyl0TyQSuVCYBUZw6wKnhG2bX5sw+
2yQwkw+gK3B5393kx6u+KLxsdmp90FQkgNE2WDOwCHYLa5AvdDLdA9lpIGkYdMHTpqcciA1AdqH2
/I1wj58bLE4gT7E6QTT/I/a7JYHQZOC6g0Xa2VEueCFDMgyKyrrr0KVYmIYlXtzkuBmh6MJlS1bc
EyAM19JoxRZ1s2jqW5+vdzFpvzLNWYOOFjhkr4amFv7Sy9voa3JHUpUK6jdcpJzqEWqa3WrrHp4r
OPzXdDPKBMYP6tNsEvK0oslwvH12MaPwOjFzZDTLp5YMzouviWmN5ptrpz+Oc8cT30hPg+PBfshN
/oEQxoTwXx358mxK1x+2TkrldnPEsmZdpsXKdFV5ya8nT6DxcnI9c2e03TeC334lZ3pW3uVGG5rD
IYrJPnlUAcNuRGCAA3Zu2eAc7JEhV9K2/1BXH08pjX3F4TMqkOxqMRXXf2rer8gH9W73U4Hk6MG+
UE7B9Ukeqx1hubUsnQw616NZk5vjAbgwetA01KjJtBfMvbxyB8qeCuTQ/0SQ50XxnhVwFOPSReWn
8BPOjJLpIzj2zxtaRsAKvecjUltFgbq5idEobiPkmQ9zZuSml/Rd31afcvImPRYiDOVEZsiCOwQj
QDTgGz/IjcgQ3cT1tQBF25mrKkd2JkQIBqheAo9dkOhsKYKKwyB/lwy8G4t3JDVdCuAhjKO6pyJc
UOOtDvRv+bbF9FsK54ORUN/moZyaBNwVjclVFI7fehDqKjjJVcSyho9HpizxEXGqNHGYK08Mt6bI
ePwplLV2aop8S0GCmTtOPVSodnhDiyYA8bK9etAdHoBKShhScLYVBdxmASYX3BLvHLc+hGUSFnJp
ee/ve/s7itzrSYAoHZgYJvFv/08M/qtGlEj4IBaIKpp1/H3EBkg2Oo20hqqqtPluwBEdzuSG25a4
bl1z+Hqbq6T/5r2Bpc9v2MRDUYaA9ocwZHbm8ZTTtwxpkz4fq/oEm+7Zp7JYEAyv5AZtYZ9qWRXg
7D/2TjOmfURpup/m1UzZACcKFDducBUpzW5j3Ov6fT2OVW58EfdGhvw+/fKLqEXDCFl3QmDYahaE
QxUF2Aw9fwTyF2vM60TI7axSHs5X1VN19QZanI8CT9azL0cY2qaOEhuL4sqWLszSzA2SCdNpZL09
oVUUgamraDAKtnqzl7yq59ML0bwmOAmhX6qJjRHEYE73I8+E1tx59xxnPnSpZWj/dMoN2YBcWd4F
jLjFSFTwtO6t+nyee24dUrREQ+pTCd1SO3UEteu8F/dV8/TtIE7S1DzeLdqv9ajRRUwhOl3yNvEr
bTS/xeQQlpeM4UzeyTBHUZd2qSfbaLT7pl6Z78uB6cufvNQ3MpUnhHSl8e1CzlMStwSe/DbXUszf
vmm71Jfz9yMoysDWd5PCQBjjbrSlVq8WXbe3J6Ej//OPNPoe51cdTSl8T0xc+/ZCWkmwsFt//A9B
fqifVxEUoqGQ34Xp0SJVPFV3nTcZgb5NCUV9x4CX0i64gbZZfzAtDjwomvoDDCougBXi24a7ABob
Net49Z+LHV6lZthA9m5OthrBgg32O9l2dhMqwS1xI0q8DAEtWMPH/mdAn6cXcF0Hn2ExyP8SK3t0
rtaa03YerwzHGIROh81fs05ipmdPXV2urNqpBD6d5I1Ka492E7oneTZGXNitg9JztOeEj+vhrLLE
tbAI7E6neT122iM93iR6ah9aT6HFaJvPqhNDNxczy0V+tXHbHJ7wA1QkSt/zb17VIFRdlVP9+M6Q
XpGqMj/JtvobnkooAnBxH7TcHfZ7Uis8qZGtZqOQ+3jJQCeemHCtiCgTZlUvvm67YZZBUB4bgBhs
yhdN6810B9p6O19GaQrbMv8AjmJ6+iacW++SiB+LCPPRwJi0s+psMqy+OX6TinrTA+NuF2c9ajDH
OeVdmNMHpjdXr6Jn4hnBu4hmZRbKmUg+X19Ig1H68EaAYoUH5J4gXWFooDgcxB/Tpm+DdgMpJhyn
QiKwSSr7z11obTFk1lh5bQgb/8AyANueT15iUWVXx2IX/IX9jgs2Urdn7WZgtpPH/t9E7f8H5pCo
dJNKK5M0hi3Wn5onJRVkFTsH6fRtyugBCsUAWxcx5HMQt3FUb3wF4WcBucrYIEFbXE6IXhcmIOQe
vlLbTUnVmcqeZ2rgkXokv4ZHyNnovh2t0QZqwCx2TvtdJ2pNlMAZEgv2/XqcbDkQVd8FlbxjuEeT
znIuLO2hi34rq3gZb5qzIDZiVkS4+gkbbZ4HJsOrN+Qc9P0f3FX5l9mcRGBALy3ku7Gma2u4toEj
16JJeefdwk2P+vECE+rPeQZeqabXXoO7hcyqe0sASpySNPSG/CNB+03OPBcnSf7n68INwLmiQJWF
nwZmiB2RWxoJr1ocTpVys81tTFXH1asScSt73ybQRAdovRrDy6fCYr9wcbTdbjCbwM7MkMDJXtey
0QC0tyWuZfNRcj8JJZRuFlwZ9918KSVNk21NL96XdJ5HY+qekeS0/rEhFOxb8QV+4TVZPoVPafVS
NwFo/rvHFBScWOjsVuJZ7TQvbMQduhRh5cH7FU6X29NYFf79QRpFTJU+zSlnQHgF2qcPAHvMCDDQ
BvWKqr8BSgSWQxo4zrnz/TMCa//g08I0XtHL22dmqRqD2a0fs7JVCdL2j6mZ7a2H/Ewb4eAjUCjV
jU7luZwa2chilyBfwiWMdA4s8ZE8GzqaKEETq5zMzs4OqUcxHwMdyYU8oCc1QZaYu/9v7560UH8x
VKFDUtdTLzBakgzbDhehrscFgiqodMeM4Yq4nXogllVrOcK0TI/Il+yyRZ9sMwiWdbwAvHW8zzwB
/UjwVO6HL59BpiQH/UB341r+SziqiKqcDKQElaRgOxQU52BKe3Q1SyxDJQVETRpCGR+wZh5+k+vX
JXiDkJarQn9glZ4NBqAYHIZVaGU7VOtbgOfum5oHxEGwpZgf/tpvIel0h2DT3u75Cbo8Uri1gT3k
GQY4IulmijXvDfHbGrL+LRQtVLGhfMxKhuEUoS/2asZGLoutlNJchKFeS+VFddUx1sTZ5UcciOP/
n0+jJWf8Wh3asTFEmX8kh66mj5vmhI+QXbtDtNnA6GigV+d3qKSPmxQYoBW38+ncuv6VRaWh/rR6
IBEA2fl/RRkbUyDHKVj1F3Mv/ZwBEfeaaaCK4LNMl28EtIUBAACcZvwd/rogp3suDaFE+QLyrXVZ
bOPt2w7m5OxbTd0VpVr5MpU0iOPtFuXO5d8ZG+jFyJY7MDtFYhBO0W81baFYQrupJX75dI49YCPm
4r5OkyIKtdd8BPhqH6gftzvjqbJ+iW2lhtQxU25Fox3+X6S7m3Qz9xGEQR0QqqOLkJKbgYZoziTh
Xh0irF5RWCjGzhTLyMioz0CjIxk+LtbRu4qO0PhtB2m2G3XiLbXxuQcVFv3Pp6nLyhmoxKqYaRbk
iu0mGVrmB97nrlFCitDNT8o8p6f0lM8CbNMAvM2lK01yqpJ76HxRvLXmv4M0qRcOsh9VBddqfYFc
Htm3eOH0NsClzWJU4jpYnubGll3zJqjw2kySBM3fjzWi6z3A7pKMxg8kgolP1p73s0ttDZBqCXHx
36nz1tVIwYo54OrmebkGlw72oh5vwvKKyAQAbyMW+8/iLGtvdukIHWZtZdEmSEC/oDi5zJ/GNUZz
xepavj5l053DoENnwnxREklRozRAbuFFHXPsi0OkLVXxiStF37lQz6HRabZemJPueoYrT9liNxu2
iVuyE6KjkbjBG3LSKhgkgPNHdKXHSAhlJ04TnbCQaQbsx9QMFLStzz0uP9L7BvYEcxlS3IH9b5v3
wrxHhIvtfV3XFVS2PIbB76awkbY8YB23k9uTklTCd3gCHVuDTesA9qwASowihZkFeNYUoV8PK7st
P4kbOJ4YX6n1LzDidM+1PrW9VCKzSOEhx4zDsYABzMG92ndTbSqTbyIopCcY+01BFJlXbkWL/jvS
4uyC705tg+0L0PB7DiYnV/mW0mE8BgXZWIz6AKZvXUmPgkVIbk+PGx443WJQ1XwxKa4xnB/U8Rm9
YX3yFo+Kx5D2ckTBOF/4F30R61Wai9oXKOIFcidg+MTipvVZEIShjX5/bpGd8fIywh21g08cq7eC
qKnuNQXxowW+ttVzEbOPbRd1Jp8oqfB/hoArCyhZ+vO/JHm8Kq/LxpuS59LRBbWad5kUEQVLXgEr
I2FKFIM+AZ+o9MP0P5EXwilsMgPvNA6K9vkOZH5gZRdUuBQCKEAswngR7dfsz8irE3QNFntId8LV
r7loH/g2xplJoAFFhAsG2eHxsHwtk6AqOGR16ej/Liss5Zsll/C23TlPsQy//shzXReqlfPzzcBX
s5+majJEvqZF6qyzSBouANcJjKkLhR9BYDT+R8ahqG3MIbkbB3JqOhMGx+ZBcDAr5v9AXWiM0k+K
Vjqh3vB/JE3JdH37DP4IFnOotEVhZP5Wa3hWfr/Q4JFX67ESyQaFP4zdC426rrgC/yCVUfJn3HKc
dn1BW0PQg/+WciZaqkP4xR4exOfZED+LUG0/Cosp9IVWfTNzZiV7TcURwCtOpwqJkFDRvFx5ddJb
LT7ec4n0SOtPFmcXiWw5C0xvOFZMhZhkIq44S07tYw6/l4gPf699oAM+fnfIEQ6iNnPG3X/XgtNZ
CnPuSjNzqZ3JNUHXLdrzXycbSlOPO6Jbh2bpxqvwCXeKRDWf5tp3tLEEToloMzkAdpGpbHaNangq
BGatz8Sj9AwVaU4PVVd/LPqFGv52zXo1oPQqqz4tFPqoZS3i8e6RiL2zCCKXjECLGS+JOri5D46t
sBExz9lU6rxzbMCwd95+pprDL403BW1Rspfze6141ealQ9962POMqZENFWnfb2V/deu027O8A0BI
8EsW8ukyM1UEN7/SyVjeEBAFAvt8dC6zaUTxwGCkNBDtKurFcilDXf5Cxy2CQFrYQ7UIpnXi6MKB
dXUbrtoRSBqspOq39tz0ah8qEuQDQN2Y8O1s40d7rVXUaQST3WXDseICkry9SQi5PYnWzS8OPCib
Tq3IS8xFIhTGiTpPZEO+i4C++zLZFMV4PbiRCQVogPrUuFVUaxSwzCC1053ic9wKdNEP1raior2Z
Cza8HJI6S90zsUdfDKum8x20ScIBWA8heqJJJUWqhirvi02VHMXdiKc7qO/G2Mfy6U1wKO1GINyO
luQVTlNYXI4OOQjk6LG3hO50DOkzc/P75HBZJZ0YkbpjKRTpPqnlB8mE6LvaFp6pyea1y1QmFf9f
yjQXxf8f2nnv08jKKSff3tfGmso6//0IR8PGU7YQq82XArQcorF9u8tFwfTKzx0ZPoDj47i3PqvG
GuLieAN76hJvXniA7e29r/5B0Cj5ygm1dH0axIfv9sbeZm6kZARtYkxgblebI37ssN6D6N2Ayhd8
O2jqCYyeHIcgquQD0ePu8BtJ42jgaVHlyfyc9NVuaUYmlIU+mCXP1Od+p4KylhsJPaufOdkFrkCW
APgy09zOyTG2HDXaNSBYFqfLUlIYBNvPPitr1SAjKejKEujTuMJW845gLui4svbjhCMKPWYPT8r9
cda+HYN/y5zJbeU3CRMnnV0Ga6HWjph3KCTfy+gw69CB6g4C4mm2OchY0GUGq7D7YypCNI3O8YoT
3WXfI+2GMTDCFZw2WdtEZfKV0GrTqKSyJlRtzZQm7QEl7U4sr9HBmC5TXaofphtlt1981aPpB2u/
1ld2aNBuQeZE7MgGd5Ub62gPuWZ0W/3fwn44hPdI7D+RMcucuPnJ4aRUoc55btsPmmjc1B9J1cuZ
ytbVJU1rUu8ld8sa2w7qjEeV6FENJVsN9w1YUtDspb3qZogcL/8giWBAq+SKVc0wS86nnydMYJeB
X3xZGgkqPz7AtZ/2ARj8a3ayhZVQqHY6lK0ocKjRiBmRiRf+UYaXGg71VE0HPPMBYFzcmDoUPed4
plB0ZBpK3kdE1J1qzQoQm8Kj/5V+hN8pxHweAgM8vZVE6R8Xn+mbSSq24vGjLeJX1SdoKWMs4QL8
L7/BanJWU8feT28px6uXLCT1ZIB6eZVHm7nK7+r7P4us5tTUfB5Gere9K1LcvOxmv8xVxxXM8x+r
ENa2hU4AveQ5V9x/Q1nb9M74RWPiZ06Wf9zVzBLYsxvtrhQqHYG1PDMOPNIghHwWHR6M+vhsouE8
Oqo2KeXg2BXGUOm6xVdKwZhgLsvAePJYATM5cybHrkTwAJgtTGQJ8SHYrgFA1pIpY7kDO5mfUXYl
JS4e813PyWmUeAFHwy8oXNf6fZ1VNFZOgiE3d///kmMFx2mlrBg7eE5bp+83BwKnlQXwv3xFH9ML
Q5EWogeUL4s2vqd0GVn6JHril+72y0qC6sLuXyUTV0vFLgDmfmx6TilQu5nNAFHEZmvYGub6lAV8
tzFyxnVc7GNHtwFntgrlnWKMP3AMy9oSGWQHKvFcIM/1wlLMmD93JOhAmhUWCWQRkQ3f4esjl0zu
orONiXtRat1JLlWaX5SODDvzWnQyORV3+ewzpo9ZddycRgefu45J1QYy9U8NxpJHDFrYcsMNFKWC
qNs7owD/kZU6LF5Z1xNhy9e5EfeVVtrboDRG/FVDEEsb30+bzxNywHeQZgkoy2nXjBCMTtTedZj8
VMNwhRkOu7+yrFRks6At+ZXGh7TiXmsq7bxKmpJTQKlDz+x0WcGvdwt2qlQ9EyQ6drLUYHqefxby
MAEBQQeoJeuXT6Lm2LZF875WufU8qT5Op4pRefmw62a+9bnNmQOB7DsQFfltnQrARciHmJZ8WL31
t2Gwvl0r5B7YdhIjSm8frG4sanU0ZsFJkhPZ0UY2bFi7Gu0T9BOxv0toU1k5EJbhzcA/SAwnrgV6
CM+KAuW2ip1OOwd91xWkcnzpVwfg9xYnwCw3Sfm1mS+oYydPVq++lG08To5ntxCKG5TJVlnkt5Tv
dZJ/kLXqGWlCLaeRZ8HVbiAklPuUf/STCOmyWs+3JEHFV7vyuAT7lqKROCoV/JiIanSXRNyumLh8
jFgahL6hx21kXNF8rs8R9r6SrmcAHHXaDuiNniJwVISsUr9i1so4TmfWgThU6jBfIP4B6vgpbUPB
Uo1nghjBIsgFKvhY3RckzvpBFadZMeZ9CCmp6yqKFMIvFMEJHfEoueeqAsKpjt8EmumWB6IezqKu
zdoh6T3Ko9/asV0r7vkDOB9OybH/n1KKXpFaM+WB0U8SlAPhVNsX+UDk89kqsj620LTvC2MgFJPO
YKxb2nhbebLSO8uljJLoy/ETkYg5fNVcBUAQbt1uqt08TqnDDejnm0rdAMcKZILlL5khIu4K42fF
LnLCSVCWLyF88M6r/PcIwuqfmYiMxaKzE0ViFr4wfa4pwL/eYNGyfhMPqigmt74hulhP9FEKB7MR
xasKQN8Lw55E95tIU8lYxFugY0jmPb/rsrqKl1QR1CMhmw6dQPuMk5icxn4ggW/D7gBFkYRoGlvk
ce11HRs4d9tKgP0hELIaiMY8GpZLWSorZJPhWfLVZjO0Kbe2xAqoOXJtyutHEUIen5ixBgWwP4+Z
ua/uoe0E9axw+VRfqgiCHxwCxlAulbPeYZkSNmkeAEBP+nRH+fxjNZSt/dKBoQkwYbBQQhwFPUYS
B5IdjFogptpAEkuJ7+W9L6Hf2m3uLRFGhaHj2EDPsC1ZsDNpT0aBJJ/RhLCKeVFr019J/Dj/kQ7w
MiFmyLC2xkxlmVfTQgoYny+H5EbTr0oldqXpNjquP88MoOACJrFC38PRbNJBqq9cDsXkrxoDJ60l
XM7o3DkzGhJRgUU5/+tBYMFpv3QLdQBfqTgGAO+bk/KCuyFLLFYI4CC3OUglSOSKTC5axvO71TfH
P3x5FiTFKDiVh8X3zqbEW/fdfRp/rlMI/kwrXZlDe8h/+O1HtkrVWKmxnH3b7t7QcNTbbpCrtSR3
jbGG8CIxMtYMNbCb0e5LxXUl5pEgtx1y/7ly6mlVuiKdI2VpIDqNevIqP/aHehxeqXBjYf/px3C+
+R4bQO3KF6mTuFkYQUvcPDJD4YdxeA/e4Ba343FFmAs80xrNz2kpikAzapF9GIUgSl0z8PqQ3yiQ
kZfMy4SG5Sg2ko8vgILW+WRmOkuBJtGkZG3kjhwqJHmC8a5Bds0vrHEP39VYPoBpdwxo9JyVbH2R
GARECDhpNyySx6lLx7c8nYuIHp2EVHOEDqUYsavrZk8W7meupXfbwfsbwHislhZnnCV+eUNsj/+C
6KGC4L4eff2cLwEMCP26sV+Jh0tP9CFXIU4+O1Jw7uCVL49fNaYeYusfg7vqEFkBqOVEp3Sd4oEs
s1QC2b0MoOe9B9o0497ePq7P1z3XQv/eZlmY6ATzGbOqgDfTf1A6x2lMzEPymu9Ospua6CpWqz4H
LsZ97jWOckpUsZ0ymK34GADv2R8yTIXViSviCPwYalMqeDpPzf/ePRpef0U+rChkcGBb4QvnukXF
n1r/FQpMhViV0auybs5GcNNAE8TqWqxhIHXC7dOGQob+otU1bVsZCkfQoPZz++IgHuqp+oMx2AYD
zGRZTfevqqmn7b4sAM7EcUpian+bOxWFxn+p3KFy95sl0Jm/zR9FC78/J7mb/0bmrQks9QkKoPK3
PUxOqzMx+e756+eIi4sZE3b7o4XfXdjaYWAmAd5j7KqB10OLRxjPZqDAy3ZU++OBz/JfB30ls4Bu
/LGre8q/ScbrK5vI7udLbwbsNZJ7TUG0xzf+eWI2SB6fBQiJu+hLS2bAG+PB6gQ2ntPJL5sqz1fp
MhuxUqouQvTeFeCfYJDdHXRQpaPt2tyfop9J7yd92n6sxhmxGOL/wTKgn6D7WUDJbfa5IKMf8CMZ
Xq9cX7g+wZI2yuD1qnKb14nbfNw6rODTOB7m8ZNz2HlF8O2jUvk0i/jnevO40pePC0ELfvITgMTN
vYiOA4Lv7kwy9Yr2oggMyuEd3juPOy2SZwMT4CheMGP+hHLHhamqahKobAhQ+BIbvk/MxjsqP+DT
74J1qIm955DQRdunLQ2E5vMHMhhf6+fkDVi8NKEKhAZQWxrpL5LbHdCRl4Mh4aKnp1WehNKWlr/A
m6MLZOeTAXEquTqk3tuDoxF+0l+/i+m3eAPmjLbEi512iGrUFMw1sy24ek0SV9ZkxkhqZZi0AapA
OtKFjFOkAXQmlL4Wmm1uLCCJpMxxgapYTbBa5qVpl/F4GgWb29yDz30WQjhLwRiuZ30Q3nPJDTIl
RxQneJ6/ZdVkTF74FPTNfg+6r6I7VfYyq36wDFsc6a75DVzJEYuEECHu2ZPORGCft7EiPKU1YZSY
WXmkoI3gVXykgoob+V97ElU2Yxui1V4vlgU3DJufYULE71T5dUf6jJYRMCISrfjXpmMJJZvwVU2i
xCMSM4hY9cULMb8tXuawEKr4E1Do3VEJsKGVz2WK1gtPQ85fMQUJdCZwwxErvaCHxlPbNvSapCev
re+qHzRarK3mPR43PKZQU8MI7IjPYVuewKeXhNSxX2hm6R1B5cyF2ahWj94Cyd/GAixYrkgoFsCV
MVMntUxq7kfNB0wNFFAxt9ukW0FN5Ko7w3xoE/0glb0ypRpIZEB6cb4wBtGzXgooRp+iCR7NqkTk
dExxzEeA+AD3xognQlTdAv+/Suc+Hn5sxKoTOGyln8lgBrvVDCkR09fW+8nwe3jnlAYm8QLsCnWn
o3Js0IxyYfpqvZvUqiYLLPKDUkP0MpuBzrzDMP5OZB7q25m5vGmmwTqxkI5sRkA8YTtCpIpFFkYB
h9p02vBNKnonZuDeb3v87930gpmZNtZsKYFsdg1mvOKqUD81DzYkBcHnTopOWL12JJeTMbjG0uhI
Sz8e6V2KLDbfpaiJlP69gRA9nOWz03awoBDa5Now2F0dm/Xog7VdVo/erTjhsE1cJPrzh8XJQ3JJ
EBLmhLfkVUme9cIVCWYN42knb+hLoo6PmKQP8gPUWTLmoUjKNGl36u0TPHR9nnpygi8fRlghZ381
5wYRGkRSbfyJC4A4Kvf/6+U0LEqlIuMa/cjfI7UgmMbfP7U//ZjLx+n9ztoN+X3hY6STkcZA9hjl
TsnAM1aM02r5BfCyQaoRDnwSXZ5G6yYj50SYn9AgqaUEuWjWxzagLQ2B1LIl7WdrJIkT/wwZ1yu+
Ncl2TcXgy+Ke9EJjRcVG3IVzwCz/2m/iVX0fpsZlZY3jMPcCpzTOFuKUO2QLGjU2VXo0G7dgYaHK
n/YyIWIGj5f13yqwVziQ6fthKBjL3SnnMPYoiTFT/vpvzb9/VjAqpWlYDQflT3+p6GGdZbGPqAQW
5n2hm+i0oE4Sv3m5bzihq6VvrFBHR3YxAp6oec17xT57hQrs4ogk1tQKvIuveLFkgTueHMm5QPaU
tGKqKkjY0P+vra1auMefSDurug/XHkVt98zCkJNPkE2MziJZLy5BJzU218b5Ckbw4M2kBaOU5B9n
iYMSl/PZUOli44yToZGB9xbDZa9hCriebORNF9F0k6f7whCDcNoW4ZAFMZc/8qtbSFXk02xcETEF
y4og70qAW1GVpJF5G9H25cXyWE1i7g6EhyNOA0nQTBvJgtvJIey67E6UbNRtgpwjLwlKctU6i1Sk
FEn4wJReUS8mrWpYkjTIyQRx+iM2bl2XkkV/XPUHEgw1CSHZJdmpHhV4qgzVbFC5OBZfXs9nQsMk
5p0qTIcJPYQ3w3F5PpypCDdsbJnDC/s++JDTOfFeUx/M/7TZGZF3GHMsqTARYMRJ0PyZoBnacMlx
PSKfqTT0lXzWTYTuZ1vbZPtP/Kdogzi6dfVgU/y7WCVNXUbYDlmVotpHV/nT5oLrLXEoDVPgV/nn
xbiKqIS/fBbzkCjFne7GKkZV2KdAoBfqxyJR5FsboCZOSYW5hTHljxnDI65O0B5jcYnQmeZ9I71j
Dgme3oRMKN2yn8sFwhIUIxLSNKdGseJkVRDuBnlBhp0aryXduKPSR90MquOQdhdwL/HitLV7+eE7
Ek0CT1BjPFU8Dz8SiKCz36qSZBumEEjS+GacRKJiKUrUSUijODl02ak0JxaiiZtrZwZQVOwfDraZ
QGs1FWLO7AD5XOoL/nlMGQdrO50LI8m53csXvfyZ7LKBnRnZ0KxvzXG8SGxgXx/9FRIaGXNBIGhc
Ft3zEdxT93K+IHaOzu1eA1RGZUL6ISp2J2N8AOhYL/3rlCSEyt8P+RKCkHefNkk2LPdEdNPDw3Me
+UC4BfZ1OQKFxKVAxemZ9OB/xYhG33WlPZzwJ8N0iAkX8eMs713IfK0PLtOpH2Tx45WfdaXdDCRG
Z0GyIWuTBsrH2gNWpsEb3+dBr7msxI75LI0seNhMv+iz9PE90UvlQBBywcxS/3i6f6HIbNFWa1sK
2FpuqdZMNKPrkkqq8XTUKuXxTAsAeG0kYvpXV8C0S7+YOejrdTb05dHyDh0P6op5ctUuGat77kmh
dbl7w51bitAobwcefKtfGTI8UifxCx0nFcNYbVr1W4pS370jwUWQc93WGtOafJ0ZWj32Zu55dJ8Q
aaU7HZlFYNt0T8EOVHd0q8qSjACaUdZndpEEp5VMNJVY5EwqMecrhqas90QCIpU8esHwP0HxYPTr
J7Pi7JU7wWBnJb1Zl+iEv62k9fk+fvc919bDY/tLF7t68I/gHnzkqizPXEDdP0izfjRS9G44ByvV
R3PUGqagwRa+9b0g3v93sP8MI2v1yoRFqiXk06ZGNXsmFvhnk5mYI9WTWVytZFBKd39oEj6aIqCC
Iv0cLf0fcikDA340YQjchjQeWe/cSqYgTGSv2PFF7rGNRvHruAeKJqkLPGmipmYfAUgCCjYe8t6F
H0QvkV7b1z+dgZD7c5i+QP+nwc5BW6ooYwT+YOQfSPumxFOVGuZzSOAHzpTP0Ue0I3Tr8pGsdNY6
vyb9PsSdhvZZ669/ND10sjT3Lps9biY/2rqC9rPqeQAl08X+Nce9+Sg27m084LwXtCUqYPzGmE8r
jbPdL7QZX9MHK/NwuS2i2SVJoKPYIetnz52UX4OJjJmsZJco73DhCtmd8lM4XwwK7TTgtySv7g/U
786+Ig40CSCuHpYW1f+M31Zyv8CJgfBRBCvdPw2zfQTvFtjciKf+ThrzxVGVZkGOm5+rBsi7pCyW
nwYoYphb4ColpxNr+0oRA4htHC2ymhE8f7flCFzGb88OjMDVgaclx0sszE400Y4r4YKCIN0c+vo3
pcD3SJwievhUTwDM5ssvVeihPj/2tlu7V+0UrLt3SMA3KrpaZlYyhHdxDVJR2sQchQfqO5LSEFEr
jIEh843HrnGzKbLs1WV82e+SpiGi3SbKvqXUB4EaM4weTpVMga350coQLHYb1N1Va8JDqC/G5njS
YG4f9WXFOHtWGDs4QBNslI0lK14DjYzC8enAj7i+OR/lsK0+qYP1EhjEDeqxZzvUuDB1dDSgl32p
xkaQlbOrfKYRvbGYXzF+FCrJJyqqxm7Z/5fDrZI85hndFH7byLGSyU5iqNhtaFpmkThYru4bF4pw
6ER+lY+OncvICacNBeIqoqtsVKw1KL7O+PDj6G64dWlr1KbfqyLhf0196sabNJ9Y6zEP7ZASBb8t
ZgTJRa4ck7DwfyT0fdeM5gp/3bBesbB+nCtQhC4RzWvB5MYU9P09INXTHgSAdO1jD4kfKGdQ3JxA
lp9xYe+swdxzt49l+u0B+kJdgCvVlJ4s/vr3F6omzIacQ/6PAqLyJowijCenSMx18FfeYlmguCE6
8jGNdcrVdEoNsfbkava4KtTIElqgVOOtIdTeIio48rh2Tz1nVlqZ6HNOWGrjt94bBwJ1ZvTRgwat
dUe16XIO/Zm4Adkx3AsUkGgYz5TrY8Ddv+qM7o9Ot5bEJJzaiNpJU2AAL43foUG4jQRhmQrRz41U
IlHwUW6tc+IkaK4Oo3ghRkgajMwe/MoblEMpTzMia0Aab0sGShqE+TVE0jMB24knLXdgcYDCisv5
IHwLTGDwUVcwUajU6bl38z6V/KqG53hdD8T13cBjLoR8E1NFbquqxAxP6ALwFjv5NaJNhbvJ1fAz
YULVKRhZyOqxfAph+tgAcxiI5DyNGmtUTTT7L07pdJa8WWfUR2BjtEJU3w8Y88+jFfW4VxaLwtAP
5Ark6DSS9odIy/EmEB8kzfKNuBrVEkufeubsDKdhPwEFwNV6pudJfB2zwkVae82DP65tFULL9V++
eI21kS269Beh1SReAGASKlpZETlbyx3EuusM/MkeTxNpn+qkPvGcXPY7Ple1RQ1TW1UKFBVLmyIz
SZ6+URAd/RxN4b22qspBz/GAZF0tHMvGqMDPhAYfjnFi5tS+hPbb0MaCJX79mrDwXiN8JYcjba5t
4ua20wD7EA1kzZXymOFhNuBjm/KXYJM9WcwpS8O9naqDEBTceXRuCvrGAMUcaE2PsWvPYC3v71dI
ylNuG24t1plbGhN7gDGBtQInMdhBXTYJRklRcEHAMSWrXli3DcRWZ8VgPD1ljEkNn14fmRMDEXa0
lBX3a3oQOhdQbWp2q2kMLm8LL5nbEkdTfJMCnRurBeB7x18X7OyEXd4nEnS93G7/6veSvqmwG9PC
ggvWIi0Zj2jKPRnDb1M/PfywFpGAZqRe3U6qWH6aT4O0E4uT5BCvIl3VE9P7sHj753VOc/QEZ3wR
MC5V7HsqL9YzgLzHr3lx4hE/V5gZiBSO7GTdG1R7z9jy44lonSZGJO29WpUWvwQcpWovfc82FtFN
aEsUwrjqUHEPjXOL4K3tv+tpT7/3+gBanCEgTYRTalRnKSQrGEN2Llex9m+ihevonRF0YNXbU31K
9OXyjtTtNgg4Z2HphtW84tQfP0BBBF1L3zlJLxeapppRByF/kdZjttMc0YRCdPELMACgfAm+wPUd
3c2Hq2+eY4yR8LXy2OylemtYKM+JGmw6nrzLp3VyJ61ojhl6xGv185xxyq4qNKujzDCcGx4vmEIk
S2xLC7Qa9JH2AkmonTmuN1qD9rixGTYNA1+1XgSZR1o9BQ/iR8RAYx/9Wp7+IbZjESRxM5Rv5NFA
OhpdZnUFxtiagNwfp6XuYQnIex9zmnPsmTGP5D2NKsu0vcbgR/t/RGQAB+u1DhbGfKEWHPARal2k
/+b+GrKP/+kXPoY2rphwwbnklk+7ulUhoKIvxMLD4BGDN9pkvKDXNlC/+rK1GrZOaPl1tZ6PgMR3
8mVFdnft7rRitxEQpDCgisP9WpxHbY73tsWuR9KryKcP1sflp8/48JmmJ2BRwY215bFDMn2CI7LX
XuctF/mVuefWh1MZANO5KNIU/3y5w+ZHLRgMreQx4tABrE0ymelvi6RrfbYnZbBq95LOa2LX75gb
rUqlZ8ThWZ+96cGCaClaoM3eShiLWM/XGQLqrI4r2N4QTW/IFKooK5Uzzj3gKC33jKNIkWP7beMm
qzwS1v4/DujkLFpPwNhW399ixmQgSdvu9vmdXiucBYMRXXY6DVnfS4338qP34UmvSs6xZ5S4mQog
OyBZsU3GddnastTjl16R9+UcnLsb57lPOHE8D+TOjXVYQrtpafE2nMZVc82/yfv+t+hs6Kz1V3SB
jr0S1unzTfEkRZ2SzVpcyUV3pIp5Amezy6H8R9EIILDZ3OYgPyokzlPXV/Qv5tBTk5JKsl4lpSH0
VpzAMPfXeaT6+3iVch3mNkZDVmmOom1o6dMYsSsMHwjNYfQh+e+yG9ryoxO1mae/szBUAf0FMYrh
eDAfQeVuMcl8bG0bbPqya7nY+yBoflqAZfh85dz+dRqdxy0dWZ5RyXR22l7di3m+Ayl6esSWCkIl
YQsr4hqzpVhhk9Ya6kfImYzBYR5l8w3VuUvLBM+lgSTueg+s/dz++uVpYy58l3fMyNSEjhKhOhwz
LMEiGvjnxzfStRqgeWKceOm3XZHvM3KNH/S3H3oWu1EfekQx74DoBlmnUX0Djemcs8ThWCi+uIfC
jaoB83/cQouNaxWUFOLM/gFxtEEbzQzBkzNnAgn6gNrzdpk26yJb8rRTIGJND5cCUsS0Jq0qIe0n
kgkum//QP460isOQFFIdiVYpELBff1S/VScMaabZMaDJVQIHQJfOrGtdUjvv8/bwqS5FAuv3V7/h
tDSCY29/6imDY8fyOaBVFylj8aP9i5elNK5WBT83oaJ7pIwNFbe+OpOBfnlwcSDmgRIyLQ+y/6Yp
hBHNQhN9ALd/SJIzyPxrtT4MYnYdpS4LoshlxrXupxd7qV6jtwQ8glH7gGMYGqGHqtsoNlf+aO9M
u6O/3ygLhMMPZysphtd6UZoR16t+KU0kPi5/skoe23fby2V5XtyMTUnnLJW0zxBIbS45eIn9ROGc
ZDX8FgO3G7kPY5GNfEIA1pKHODkf/EyoPoaZ3YeMMCODUjMZ3jFz/G5vob1me7KllviOTXGBaOEq
SBuJiAm45v40NdbSZV3904mnNv3yF/V+eIEQEHVfqBGywE9I/51yNery7DMsdHUXFagIvNRHhl+b
0ZRRrJp3pDI5Ilx0r9/I8iX1rc3Hh+8Z1bxd7kj1OwDsTXaIY8RmpykNsSw7sQLH0Yb/Eaf4STDG
jXf/a4R9SXzSlML9V57yG3RLc9lnchkXi2JaEYae6k8u9FK0r68atbAfqVyBeehMwLrWsdCQlCaW
MdqIhISQ9n6TGddNRRZC8JwT7XAE6Pw0fWolVsomlBuuT10ZLIBVTq8aLgGP7alinvAR+nxcmdFl
9tMpmIGS1Tf0BaoORb1ITDhVzteIBn7PyhW+7yzb5p6sk5hMSswnOsq4E1V5xsCRI59R5FtlmL68
6elM2iGbK0mToDmMNqJZRHbp/zhGDxVWtTgRYSyr1ZJZXyM6rUhCkizCmg39YWb2PyO7e++E7Zss
ctSz3+tenKGtarSbYN9d9NHetfw9ArBo15k5dznlraX3i7l0HE4m4ItkQkOZ+wq88dI3yZ/s46yl
6LwwLqyKKRiRGfDO7CPncnlnlQCYtTj3nqXjuuDoGzqDIuaX6hNuLwHmr4Q6a+iKtLNHz9xxsYz4
mG937HjJdRrXJ3LA6+9D5Qlii8xyGy4Jo3Y9fuktmmaWVMe3NL6icuWuQcSoICBfmfIavcBMaOt6
/Dy5/AN241sgxDHYOuGMumJ8lPZHFtWX9YPpi8D0rUy3QChqpFnef1E8wsDTgFBYLz+Z0fOd21tU
leTMxJA4fw6ZWd/KfvFPE498T1/pAsZrC1rKVTTMo2KUXgznQQkkJiwZZS8SjLxP1gY6JXWp+7Tl
cvIC/vqr76LRwCxF0EHH51sHAy8dBu/y5T3NBJA6OpCm4iRFqTejF6q0HSLYuquYxAWmyXUW5+OM
i6rBUShUhmE2kt8JBMbhHtoXfECTyoZh9EFlmTRJ8KVuBdpw2FXhKAfx06i0LTVjB1aBbm8f8xU9
JOR1G43fTx79x1bxCPkr16KSXK0LL+8klx33hgPflRkuot2Jzb2IuB+mQd8LcLzPIkwL/0T9yBeG
QVoxxqYpBaQSW4glGlzEfhZCELdivQHP5fhpBsOPM76wRDf5Vf9B19MCtubUgf0CxnJjrgfrDtMn
U5HFnWc7QYnlY3Gl8og8xib6rd9Jqm607LsQI6wXwVKXe/W5r/y1qCKvlvHzeGOB4K+CvdfPAIZl
yd6SEozLpvg/RTQNpIekcfg+pVqJ0Q4dSMa4OmQhiqQFp71/Aeir9V42+YHTDSXvANKk/4Id7wW6
RyBFG5QF5EbcISCD02GcH84OHpkgdWp88AERnhSpmyCrxGHGawW2ZvayBhEdk3B7JhEq7ILlRH2A
oJlFD9+mPHuYu86nZ4NcATtGGlPgbm8YbwgZqcvZ3Xpy78nJ7r5YjTst+pwCmP+ywygITW02eAbS
gfDI9yTyYQOzlJTfrLhWiRXM1Qi8hn66L6FY727hNjI2IcKoWOcYJkeGU0FILZa87UO8AVwlnC5n
Fld1ne9+JbQOaqvS3RQ6Pnpe3JnV7kVJeIFNDhvtHwCOzo0Spkb31IICBLVKiLsbgdGF2BggiAnq
rDsVPCq80yWfVKfa4aW2zWXWItHZ5jN0HH75EivBUrzjzkOJFswFc41aagGVcSMf8/6FCwWYnfhY
xq0IZ98aUnC549cC9BgqGoUceFxgct+QgeMtBsEIN97fT7UfZPpD9gNjA+WofPc9cxMa8X3Oo2aY
F+CHV+G/HfHGj8VsZVPr5Gn9hqSaE/N1R4cJdEi1rU5zSDnM466YUZyJTTlwy09E5f87enonRe04
VIMRIe0Vb5yph90Y1H6LpqwWRFiXTuBTzRVkfo3Fe2WYBx7Ia/Z7igKLSDZfHmdYbN4Ynrq4Nv0n
S8mlnCVibUtYFIRprqwDVBH2Kv6W1OH2bztzynJM7NdLGwntspRWUv344wXkFX4HihmEt8H3ZOEJ
V0ajvNQOzzfiE3M78hLvYjHUBNEXWLMyUMSkR82p+KxPuvXvJuYNOr5qe/TmTWY+TJPJyqKweqda
JOUZMvTpIJItiCPJ51n60yhdO/d0mDJwUaLkI+hzfApQW3U7e9KJE/Fg06093ZiyZWBjuOlABgug
c32DerTf4pLnmIlPpaEoTjdc1Cm4OSny+C4FdQHWbm8Ntq1wzhFROmP4UZx+x3UINpbdoEk5ttuP
zjtrEvE7C/lVT48e/7ibzu6WeLhRIACpXbtKpetcCIKgERK5SBQDb7/JXbhzI+ptMMrwOs8LbBKA
t1OvMOHsu+t4WPZXgJfgw5jf2C/6ql0Fn/5erc/bN95ywMz1i/xZ90jUQJOenjgvmpuXLQhhDh8g
S/yHmc1Wnty+XvjBcsqVk7mBFyWUZjW92WGdDpaAqp6n8qjgEfQ9H8LuaMclp+OE7WVTNbx9voly
ic+BWzdVLSsI7JFMz8lDe4jaf/nuXb2dRqGY3vu1BmOgWv4TBtKNz3M28NNGkPauwnnRqnyv/AQT
3Xnz13onby76w4Dlwqg6WWAFsA493bGezU+YmpFSrIKHGyhj4PPHKkG0LbKnhs9mCwuhcarl3LC3
9cum+E5C+hWXBjmJoDqjoceeIs68tk7xuS8d8Xi81NmzJTSh7BsiWFdobmRpY8xCPXbT1T2jmSTa
T8Xws60qVI2456sBsf8He67XM3xvroYJhpD1WEih0kUzkPiPxhteYDek90oTbi1W8Cv/5Ej1Emf0
AQEIkaZH2c7pK/PymlFRNu6w4pGPrEIz1SHqDo67kugLtB8FvNfxsBXg5oeEM9tWZ2JIeHRchejB
m1jir2GtqTLKxQbH2ridhPZL1EvLqOtRvhwGnKhgbb320XDc0jOZYH5q2YR5pJBctp7PPQ2F9+cG
ZcJGtAxipc+0vmOgaMSYv9EYQ1QFJ5nlsqFFGlahxlP5O44hWD/MrxipNP2f2SeSnnvi45z1d+Vz
c523j0pHDhJA/TYN3mqgVsW18OhYtJzKd8S8mlgX4iV2aYyOgFbmeTCN7gufQyVDphxRKZWy5GTB
9+Sqh/qBfcO9PunafRzQIatnMqWtoQ8HHskFqcXuxw9ilk6WdwDnTb0CPabJTAGlIX0YdO31JDFo
PypK0SZDtxuWNTO6lEGC0TnwBp2pEEe2jBbsbUl4pxHF4QvUkIvLdVrsrTrh/B9ypcymF4LNuQb7
7xAxpRWyTL7XBdjuDj5X0OeKpYju88W6RTBiYtFClvEZvN8O1Ab4pVpVliR6E4qJ9ALjj10WZiKc
NFwKUuCbFnKvMNMdS70f/c76CdjjdhR32G5i6ZssUsnKkxbNHtQ8vcH6zduRwTu49iy0v+Ybw8N7
GDV5ZQi2XyMSvYX2WxV+RigTCGUIxRELco1N8avNRZAs5HAA1O4+2ASXnMwfaYrDe7TJEJesUTt1
E1Wn5t1revWZoDcYG2fvS/fXgiUctinO1cOoc7z2O3btNAUgICKnX2LnamJ0kO/5Rybfi3VEG9jp
lOgDhLLI5hrH4EkL9Er6sxrsfYKv0ILqPHWuGAwHPF0zzI2QNKsKMdrlShxt4cIpiTn0Kjbzb+IT
ACRjwuaD4fgfyaOyaldLV2+/sR6YU5OElpXk9Vx4v9s2kQDXplNd9l6Uw44PANHajRloVZi7SRqB
bFwOdMKIS6wfCbAuiKZBRW7XvnmUDzjOeEw7vW2YoaJxROoRp8iKC8UQaAcFoQ80QceIkamCeIjW
DjAOALkyKCZjiL0pa7QL+Bv34b8BigSfZp7nBlwI131KjbSSlFb5HD1yVQ2JAv2qsQe+r1/CbtZN
5O8a+WFyuHkE1sLckYsycSoZN/On0L+YR1EGhvDRPp0ZqH4pt1xoJRSB6jAXOgOQ2u3OgpBD0X37
MnFsXCm9uMf3Vvad2UmGyvj2eGbxrjkT1znlYn10aGlql1Pojw7+gYVS7PIpiShIGJ9ljfGX8xb8
nk4Rgc7YQBYcDblxmnehYnNSAWIdEd7zw50VLVSRivEhFIWO1MYLtdl2La/QJjwYaZCb7If9+LK4
AOJWcMB1d7MJlMAgZr03eRcNo0z5Wtw9wBNUpKyeua/byw7+X0va92WAiWDVD2rnYL3PrdWDHY5p
rHgCFytjTz8m2c2GC69qIJpirNR+ZD5RiVaRe1Lh82z2zJ5taARE+GJGbqxdOL7Kxp0kO7Ll1oN1
hLPt6leTukTeNzIaT9s34KBZIbap/xYOc8jCM+K+yBIwWndJ8lq9TJaFNTEf+CMasnxMHquDFtKk
Ki/aRWwoi9sQAyPN1CvzVJrWsqhtus45ngwDwZCuNw9tyzYb+0aSctg73qgAylS5gDCTOgNU2fEu
X27K354koO7EKZ4PDg+pXUCEI2CZ6GCTOP27QcNQfSILQ11RHcJKRCMhkBJsp2FcAAVDrZq6RIKn
xg+EYJD5nEFVBoKNPcJNszqyxa2Z5TFs3xP/MCL/jhj08FdjqpEa+aiZpPaTXAyuiojcfU+NJa3H
FIF0m53hSXpJtYN+FmkWDpRfqMoMUUzThHmcgLJn39SFoJlNNXyRkCooc4rod41Yk+mrKB1etwqt
sTSyuavZvaz0TwL3hd54dcThNCCk6clHNPKRbgxUmQooG+uWmNXIR3nuFcGoCrSPOvdn2Wx63iOe
RIeMTOQO729C7y32+Qr7CvkytMORlsaFLC/+TxMKvH/OZ+BUuMvIjYx930YeAzIwp2wvrzOuz7A+
Z0JAdtTfGSNLlY35F0Eqx19J9Du+CR5i1f9QRNfgvRuF54fmMPMhB/eYwqUfzFfRvjdGLmwS8OIV
Y91nFosICZ8giPXue+ONI3xzNAccbR3Uh8gpvtjqPBrkctgdM1LfxX6y7ZgPeQBxDUWbcBD0FLkr
7Ygr4U2XfMBGwhI5wnCOaJElwRz/f9dCzVg+NklbhVUZ2O7zLDTEOvCCvibslToLkY2LcTHA72Fh
5ztZ3iBMut/YUt1xGCVMKYaAAwL1S3wifaVnSV2BSd6pwgklz5UAVHPLryuMck7/k/N9XrEs2YPZ
vMccSiJ3t++aSCe1MUZ65jwkh+S3fGaorfzbPQy5ACSHQ8/fk0tRxdLmzlZ5IBpBQBqe1wuzpIHy
1QrOxo8sC8GNAugS7I/bRbgLU3fvWbPCGhkZ1h9oe9+XROYiZiEa/2nQX2qT88DfWl5IJi1C8h9V
eXUvgsADnTcVPj903b0g+/9/5P4MznIXMcdg7pgiWzbnvsbyH4TGhT58tQ2PteZGnnxrfU5JMCtx
2g/EIkgtm6W1liSJk13BeBaJORREOEF5ddEOW5QWSukeiGLC83KEdu6FN9xyy65Z76fD5nJ8p0Ee
a1h6w1v2Lj8whqysPjYPwxiRYVEvbH4X1ho+579CzaqXpyhWI/2i7CUF1d1/gRs0H6bl1xpoDy34
AE1EN2MuzdBydxQD/w2t/4zc1X05kOwzyM/k0V6JHeEVxobiDAVz6yVCfUowg2DHRvuD5mDiRIHz
N4Rb6x1SW/Ts+UWypKBD43FfVXS9/jEwhlm873lS4ppwdb+DRmiG+VfnNwgNl1tcbZD4OvGgPDdl
Lgr1kqpD9jq4ePaG6VicK9HyNgiYzYwNAyP86YilNRfUqlswfz/JJhAI+7/HMGDS3rnKsysc7UhQ
37I3hkm6rTJuIdxRvNHmY+n4TRKW9Lu+eCbatcCzc3bjZVEx6A/cX72uOW3zEzyMliuRs0M1ZfQb
28M+PrZMNzloLcQjKdx2Ttl7BdX+Tcg2n283pTRhstpJF7AxG9lkYKecSB3USWa/8/5amim/9q0N
hwybylcNCh2ouEFoEziGdX3UVnxAGd6iy34cwD8oxbYfuZ6AGtllotGHPEx45DwMbBmavfSpwrRi
rZwKDucbcvhdLq1HjDBsWXDYCk/iHTfdhsl9pTc+glGh/EmRx+sd/18n2KZ2FJGrXeIuE9GPKpd8
J0YrRiQ12fTwWfl68vMfwkJXHsZU/em+iI6u45LR+tcyg/M1trxbmJjh48LmvNEtPl7F4Mk5iwcf
yTQedvu6X4H0culMhzNj25Vz2+qukt+eKeGuDKVDAi4NFd4yQkBG143I+h9xbZnONTZWFAtPczdd
mLeaeIVyBcyDPjw84xmBaL9A5XrjD0N5GgeK4tm9knfsnbvTb/oqZauy2yScVXwa/16lJv94NS2+
GSI2i7EJmguiAGVvO2aeqilvu8a0/6Xb5aVb0o6EV/Mebjc/ooPKUdGqKpg3moWJmejpfgL8WZdc
2/CUXi9GLcF4h5rZTGTimItiz0NmiVt6dPnZ0dKHXb7BQvZ5RTdKLgPajGYkywBYZ75ZsDCa9Z6v
GQQ8UV4gXqrlRl8hBxe+KDJVvIlZV8chw4L+rAnbumFDdGdWbZenMzJYeNxRubZumwqzo3tBJM3K
rShVBOyqgKETGSZBRhvSlJxzk81CSk2TqswrQ6iPg1YUkyoQXxlNtdK5hiLdkdIvPAFPOZpuQpEW
3Dh4cZw+aaDDsde0U53F7gBkjzKtMR+DSNFkLWm093zM+wPbTjMR5mUNP76eUlY81XxGg2wUydTD
S+qBmjPkaTtpCwKjKQNxhtN8juo8/p4i/+odFRl8oyz9fNW7U0wMnM5M/PgHKb/GealXGMrtwhae
XBszphEbEb4iNTH8NlPnCIgh1RDzg9BcaD3UHWXk+SiaN9AohHzfd+3rhj1M2y6Ge7hfkoh9ab8k
/oFZRlOmvw+s4FLCx+5X/sIUvEMDGbfPvdCNJUfMBu1kHh4/kbkoO1A3L0u2wYXEcIwcg4SAk8U9
fuBFd79ZFhFb6BEPsL5TWikKun2Z9VA9cwSDTSg/sTFIzbV+u5YrwChbqCkATrRgmm1COYKKaJxl
Bd6epkGpZGFAVteIHMF5RH9iPt+eWzgrrqOPYR8KWK6nr4xAAivCFcLhpddnL330tO1wLgZutQod
nBKqZU3tR9qPTgZKKApsqa022MOb4Vv19dP8WaVb8Qw/sE59B2tQ+o9H0MlMY5mm1jprMI3QmhbG
BXXUPtBsf+5QcPtQeZ/VX7uHQxvTtrb+QZkDNfg1vmL44jX+v1iqwm0ioAdV+a6cb+jkipnFc9bV
eshib4pOcQMMXDfMgaNaNwOz5AkZAf/ArD+eiFp5B1jhxsDadiTPmAlrNoX7RY7QiIi4eNJw1jNs
W8rLOceArPsNXfk9Lnl74eeRFx87AR/9gRT1n3PEt99poqY2FBss55XiPfEYXw3SyYzCSbJkq+m/
AUkX2dk4a6O8puncP1zUsW5ZMYW+qTPVuPVkXABqiAnQqcrQsWeJYRdMlfVp78ZHkqqgEpLM0+nJ
JfQQQDD7qanh4YILeYNAphA9XFLMaAaX6iZYVIyueHSydDOHAtIk2Hlb7gag9r0j74ieQhIZh99u
CNgpGLAJQrFRDyYj1tLYZYC5Os/QddIJKticwRAd6tKfOQXz5VUeB9TVa95Duxn2B7d5AhJXz6xU
Q9w/Ibp0LXciDS8tHtpy8qM+IhmVdGSetNA/5VyMOjcQnaUjx9weC0bAhlOKNbjm8Mf8ueL41OrD
7z6eZiig95rqfNY6P0b48iGSYp4rpLWz6VN0U9jIZeKn9FtpcV1PKik0+1zH08hb7jOe3XRMak1B
qrYkl/c/qlgtkZpB8rca8+2G6d/g4q9kjtKKwhNhtTVM6Q1/+VHyCqPIFsacYH2GLBsgUtqCUxEw
A3Zc+eBvNEY9e3koQRhdEn9CdYLdIv/l+7zb/jw9YL24edSmJf7g1cea+MCpn+jRYfQqQ3giU1fM
sdgDQenbvVDQPODdIfjr/93o5YnCPmYj4MCu7q5T1DNhSUNm1ydoX+bs1F0geS1P9Q5AzUqmuCh0
lsq39w2Nfn7p/jSlnMlFb3i56+sfl03VlYySH/FH37G3o/3z5M3qXIowEZACPioVoNQVkkG7lMDL
1AkbZ2YpONoyrbmfUvNtQch8w9DrknMTYv5kyNfrSw+H2hHAKT0GF3H0VVX5ZgClGVB46SujV4JK
Li98ISatnURkw+LIzRCv4/E/VfacSZ3Wae63Ql1USOeFuq9P91ojWk7sY0OIR+feFTY2wGKofXkR
76SSHms1gq/D7O+sp0Y5SFpVPm9k/VN9xHpnDZMfE5TzO3LVZadSHR1eit5AADCVRC5Hs+Tsj7Qc
jVQ9q1NrEG/alGycmGm1UW+Sp3vyYiYtTqB5dF96/y7cgSGrRg5We6CwebBEviVx6NQyeZuEVQpk
NW83Tye0IQ3PEHI+n3QKUBBw115Wg20q4V5AQLEAbb4DVUooPtXTW+EcNg/NiuFv5JpNpvHWZsCX
EO9zbFdz6L8tHvPNS4PbEp8HW4f8ZqTJ2U9+cCx+pFuwMIkPlZ2y5VXyedW36F2yBbe+XG617vJw
m/4yVTsb+W6QxC9hYg/cLR1nZ7XLQx8HoU/khO/XV6CR4ZzyI9CcgXlmOceXMQ8+869H1wsoKFfR
9soU+SAvfwUo0pilCF5PprgjFDKecXZqWSA9DqjD67bxJj0/1XpCy5aT9XliLfyx7K+aZzVvSbJf
JdZl2oS6G1qs6rKHki9DMa2DfHQlmMa6r1up7DXT2DmdAGK24FoPxrFC+I/emvXPiJjGx2lqNkC1
5veiVXhy9q8/6z5qGHpLMAmkfbmmBQfMiKhlL7+eNEDiuSuHVvnbwxlCcunlCYR2/gDnrFmxum0X
P7Daj61/1CWIKl8bOjTXgJvXTY5Vy7NL56QpBNt3XursOzxRju+1lp4rWuk71m9lIQzBfWAuGM+j
7q8kmTTZ8/bWihU3gZOzMnq/7enPZKZoCZSuaWWINxfHXjJHwJx7y5wbKyHT6Psri/k1aApqE+Vg
PdJU9Q69OwZLX0Uge67NXbWVlDgOSkCvk6PcGFU9WuvvK65yO1u060/YJHxGPKHrrHKMgpDHcuVe
+iVo2gPrfJxOcLIY9/qNdYmjxEWHSDyr23qxRCF1OI+WsSTyORjPPFrsK3L7Ty2+8cATnKeDhrgd
M5alNi5ZhDlcmROuRMM4zUEgp+sDKa3PP2fPcoDhvHC/Cr64vFRAa/Ky0pjzrOY9WJhN+6JSAZKq
BIZWxTchW+mvHRiXXjQnF4jOjva68WQUmNa5XEdluFpzEkzp4qL4rltUTSsdXE5CWjQrUR2F5wHq
pubxVLMqRSVA3ZVLjyqoos1184VyBQJy9XI5Q3h3qXTFS4+J/a3kEw/TrwT/0RSyyE+BBXCb2Xbr
tP+1jjizyiJH30qYC0/r92Q3bQBKSzW4nNpqBbcyAO+AgoYv+kjCZHRPncb/3BAYTatOlIparFlK
11zEAeI9nRQLbrN5Lx9P2FRpV1QFITQIfSHpGaHzFpW4RnX3PXkgULTyKKdESIBbCh0BJ32hCksd
redCLZMuZvweCP95hy8BZCn3vQf+2azXkMs8ffgS1FNjsh22YFOfCjwM4LwlHGu50F3GG1JlTdYd
iFnEo+Mll7j9ibL/5AZD4hP5Uk7pGWLmlxQylvyRAoL7W6+ZSXX0wsjUZJa/K7BaxN5LY0FDw3+B
LqxBtl1HCEHZD49d49Sy0IAwwmQklZhY0osHF7lzakRhVzzQz5IMPHU7LlK9VB/Q/Xva7WA+AjQp
zzXfTCkLTKAGJyhvKogwrnTzlJYSR+4ctCNjDDEA0QQ+ue+s8FF6v6hdW8M2LvEe0ClO+3HOv/v5
R60CnC6PdvoTEoRZUWKb2i0J+vGXGn+kseeosQROj/0dtxZnqWlL+sHqCRbwCHXgPWZXUR15+T0V
66Aa//SYbw9ai3RoGZER2QAMorr0LburEhoR188C1WWmJWrrUtylW6ye9slFHpqEOFTjRHTL8q00
B1vmPcqkcq+JWQ+RuAU2/rtjXNN1EYXeLcZlquVO8A/QWHFDoltShhTYo+H4+0hcku1lCkMbS4sx
amF+rZ0/k9E6ldr1VDacSi/veIMoqUqUzvPMvwtbFzFvYSNxNFUeutZcLlknddhfPA5J/BBUZz+g
LZc+9YhCU5dpvmzAIq16iqTTZbhK7yJNAPs/XGjJdMirrE2y/vDLUbuOydJQAeAetKx6m9M6Rcvl
g74iTzZhhkKGi+z9Px9+7i7kXggB0n9NTa3fa2mtfDj+nNJuX0AJi8GAiS/uaWH4TjLxIB/Gq6MJ
kS4shaLk6hj9NTUj0yoz3E1sjXZ8GjjpxFSJ7msxUX5eJs0RpbVFAp/NNYgP/OzshN3FC+vwH0vx
wx0nQQaUtvTKvnvZoIA6jIQ/2bFKIMoC7GdSIL7JvCIOaCjIhHE5nyaSOWZwpJjUOD5AOp+T0wMB
csRyBhUYyK66icjMl8ISDFMe8oyNrfbUB2b9ZKJUZIQpH2rfO7grsoEnR3NGs0YHYCvOePWk/yn3
W9ie7bu6Ap9Uk5iQEwLmdqWrJjnlk+9LMKMltzBN0ltBz3gqfocxRwJnbCn0dxZQTyq34M2Gm8bf
xEQbBu3CL7RdlVrGWLdlG5VGVLsiUeXnoBKmsg8isdqTmfmuRicJg/d7INvbFNR8ZgiQwfTDtUrL
DtE5RS8cnKe/HbIvvgZKUKYD8uUgPxhtYX4s3IaDfbOUd0n/bSFmwDCbEm2vbCbBmz03J1J3eikI
DVt3Ogrmc8ZMytJ4J5pZVwRk7OC32u1v7vlofDGkJPmNXjAtbe/bpuTVuSk8m/WoWa3oryu6kt52
9n0nzpQuSk2R2wQ4S/YmZXzQqKI+TL07B5TWK/MYVH3yHoVnMsUdTZ02v1+L4rwtODyuWI+GyG2X
3uQFyVLxj8jXXe3a+eYCRpN7NUBkmvywhiqxZ5xuMmcLMElnoxSBCA7AW9dXa0/3VeNzecH0vb+T
cntKhKIQVyB+PksSzoMvC6Y2ztuIfRSgcG53rYy+i6QTX6jvnfEyz1gPYpA1CcUzBunf3qKt5svw
pUbQoxu8nhg/3tUD5HCKlN2c7Qr3K5n2zmA1Lq7nzarG7aQjtTsn0GvmggGmYTnpnQMrzTdItJZg
2fzv5sGtvpZ8zKya47f3slVqAbwJF8+bVYC1mrUVuB0hsOAyN5fmBmiTBTwBfITudQYN2kiL2vHo
qcSdP45fgt731scjzarM2DH7sWbcdJGIGE+nLZzpK6nIZ9m+WtiY7EyBB3/I4rfNeLfl9e87txEE
VtoiO8n+Qj7lNchDN4OBpW660x/182kWR951NvEg5ktqGx1hw0vkDCGtdQ/lkab1Pv4DpJh0GjnM
NZQ3UcxlSdsAZimwK/0H+N3brVMZaYDbyddbYWVZU4HJLSJyeyHhHStca+qWnsfErvU9jcTbvelR
FC4ytEBpIBG490NneHgm2gRTB89axQW7N7gOyGPb7NbwJXSMHc+uXVw66pfQW9YFJAEuLrJf+3qi
SOtSsmf3liAOhnPQKc0NfpR27JmpmeRRauoIt6hxh3R1Moy2+JqqfaRAZrqIsiGnsvRU5zd1/q1L
JDYh7WRVJDYxoq+CVhg6OL53Q644o0BkB/gQ1Sl/1GjbLFJD7fmW7n+ARsKlvxs9YX7nOtuhTeCu
B+Ah+5rDCjfkPSj2l9EXCmYKn8RYhlQ3CfDkTUxsGOhZuapNC6kXcRgI3RbG8h4bfCkL94O4jL2S
afTBB8lbRi2Csnbg9FqSxQ1vex1dvYMDbagYyBgY6SebrQzbqb5IDvTkzce/fLBQ5qUdu0RPFVgs
/MGaHnVDtX9q3Deogx/bq5axMX4ubFCjh0WhKAqBdZtNXGLVvA2QSKfQur2IH02LVD43bjFimpr8
XPrXHjnswvvbDne3j/MYIIM3IeKnT9dylCq0oIGw/mig+KpyY90x+dHAPhXBn7u2OfUxQTY9lbV6
8khykQERNk2l8o95rTUzJiVxiVfAGsB9lckANMWpUDdSv5lQKKtQE4LK2/4ErnUh+ljR8sPHSlCz
77HduVBxSkfumd+SxpXPAVTUT5/Hne35A5rs5Ry20eZuZl2Lt9nhttalWpzHhTI8x+B3hiCJBjCp
ngBc8hCQSGhFYmpjC4goEttnY6FuLdIFQ7n1eLLWbVSEX7472Ai0dvs7JRKG7MMhje6j0oH071+6
9FCyTKGRN47HkoOHINmUDdM7dzC3VEktRFWiW3fhdLsLO6E6HMnubXHXgtuFLuZRCOooYyHwd9hE
PIDT2kuMSWLlOYBc/VaNBm/2VpPVdjD+Q6okGMUZyko7gVhGtRmjN9TSxM0wCy+XsWOPS3UszWB3
O+gMrjAmuzxn4sQE2l7qLUaog8NBjTP6WBEMUmvMZef0V7wT86HWlmfTNnNaA7Q6DqBJTgD3JAtx
Dkye6omZ4aXnn1XpY1WEB948OVOczt6sqBVsFVdvVnIt3HM718z3UGrs8X3elD2eOEeSFUrYbwsJ
7H+vj9jFVbjq+wSmsr/EQLqrAJ0SOyxjI1PcrodBVogscaAUMeuYNO7Eb5wwCOVNx8pYyw7ITyam
A+aevitqOBNHXXXUoFfKl1wM9KDZxR2xKZ+fAMSzPA/0rdNXxMv2mkCu6pYUqo9czWVB2XHrDu0g
ea7f6sXde3U7M41uWqICBLERablkVGI+jFQ9Teg1EvS4sPyPbcdi3Lm+KFU/5XjdHooOfoGgYxWR
kE9dJfinF8hXheL5HLzO0lGu8pTKye0NCpF4wWW4ra8QP7/3gTLVlz8J4nbLQLrT0A0I6nkQPSX8
Sh6J0SLqF9su6mqVKpHRIjl3oaIhHRAGRq99uEEFpj0GnoTTVYfCIJ7KlV0ZSMHCvOw/Kbn2MJFh
ZT+3u0IVQIn/EUQIQAUmRneYIRKS0tB7Yznv6uDo1cGP+W02NFP2rBSz2IhYyt2m3AtPQb7SyHQY
oOCwRVYQedLznHwBIRTOFGWe5YOHFcE2fU+8zW+oP0W41tSXDoJRgRGSYizOAe1quGqENAKvBtXy
L3TPG9v73ciD38vvOK3yYtgDjk4YhSDQfAknkG9ENNbG4w2rFS0UZS6mMYXA824DnLr8EDFbhong
HcFJUb/vJl/jANKjhekS1P8aWGrM3dk5tNaKqzgYNxcPT6tXlBs+9kbD7yErAZPpOtZIJ2hBpXyr
2Kmlce/zhWT9EhAL2v2Di7RIdxGQ1Ilibhn7Tfw94N4LLU0T2RCcGSxn7KdRhBScrlAe9pGqU3iW
2/pt/npJundBSq2AD2VmYdvry/Lh5vwWpnmL4VMWEmYDN+ncAtW7nImRNeUfY50f0nAj5alec8nn
Jw3z/LVXt73Nm5yBHagSjFdkmG06sd8SPGMKNdyZczjoJVKYc4seXOgtZnG2Z6FCfvo3hMvGf3PA
gWO8BbclF4+DIr7YKuhdxPxNJYPDuFJKgJQbtGVRbWWzcMpTGo28yZnnAdq7qcgWpx2JTdEX1w6d
niuxsr0J5RZXcMa211zD2OKH+WamDQ1zALitphKW05hsxgbw89PFLNknQB8j5KVK3Y7zotYJfGRg
bcy+Jj2HaHuwGTFq7Ipx+nvz3mEheTrnG0LHwIqZ0nzQFhrCgsxmBMEgOhLEwDMZdw1ixwL5shdm
/Pzao0d5gVHiWTAx983QWQa1i8KU9V8JsQ6Ey6pT2/gWEsZoutnpI2dqpoipHT13xR6U37wDRnr1
GueVw1TiZwRJZqzTetupPWdcM9x1hFTys5+IrhEnAvuwf5sYD1bY8KLDWv9svqWam2AzfW5aDeqO
M3tVgpakZGANMEWRiUU/wppheF3Cy3Dzs9XQzjnLjXDCo5rynMScOXRUdvFDiYNZSAfg2+oT9I5G
VHwwFSQWN8ij1lWa2K+HglP4YVRBOD35fy021ZQVOEG1ZV2IxaC+0gJhk820tgTO1Pvbo8XSHO72
LNTk7KWZ/0ckviMnH1isf9X33rVy0PKBG+bC6HlXKSrgXSfumjqE1/455wxoRtObni8gOiFF4Twi
Tl+kpT6jI5PWoLB5YEJOkQuUZ1W8LsRBNL2ow0UtBmziv8DWTA1ymKvADK7CyOAnR0DFmsMq6nu/
MesZ0xC0Ri6UNe3SrvXVG2Asmz9L5EJmXYqsmBfSMEnrJl/6O5Cqsk871fTjZHVGbHqzkVIFXvTl
naOZiF9yQdfwCY5mw8WpKC1GJdaP//GxSC2er1GIuy1z/SWGpZ3vGs4FLCCBpPpauFIYFjnUB7fr
YVRSIWyEaJAmFTyLKA2RgHMGK041NIprwc+7TxLYtuOpJ4vLqXDPb0vS3nzsI3j/riDl0KADVEsz
twYPyTwEeYM72IOqZ+g6TfZPialW9fsgcwR7Gu7m64hMLul5DSAnjE8CmhHAc2vorwcwCujqVsaE
ak4sKaf6mWmDkFfN8FIODp45aQYAioK9/ETccXGVEX2wE6ggfWqVgQPt9uKSXIVT8Xn0mUNkP2g/
bFeR4vtpC80hy+wvHIDKJNBSivSsnW6Sqc+lifV/mOFwlZ0nRVrC4ls/cBOli0h8F1DOmNeW781a
wP0/b2x3k+kWJbUrDTtPaB+7/9xdRv3OWJcCOQbfd498+uSjMYFNGMQEMehfBoH2YaJ9AEH5qrdT
mJwHIb3WPpAm+kXEZGznsz0/zJqOM7dA0VJStFxGgCN51V8t2wPjqn236HBCb8jO6PU4UP9vaDEx
+epXsr/2fYpZzyDTSSoCIc9Vink1/RU9HWpPVKZyEZajigC4UXTcc/jp1CnWPSKgqcN8GvQ7BZ5n
dsAhdIljlBIKT2OO9EcmwbrjbL0yxia8D0DbHdy/+plNJjKvkPP5WSoLsRwn212GAMT4z416nNua
1OktGPmPmWk+mesUAEf0eJBQL3nN8cZ/aA4DNtERrqAPltpqBn6Pb56QmV0BAz+A5Zgrk6ETlPRT
oG9WMa4c38XC5NV37P4r7wXybN+Wm7uju5MgDWjnBhHbMbVaiSDo9ZJ9HVSEwfFyPn4XD5cGTjEc
9W51i2EnXDV6DVcUKuxjIvSGvhudlcmzqSYgNK0yNrq0BW2tV5Ho/ACSn7sru4OUrSj/qsqxxuD7
sp/6mpnGdiaS2i3OpCt8Nv7LY0KzvyPYXxW3SqHIH009v4AMieHOk2fwwDqQT4GOfVPZ/eODwDWt
F45FjtCkOBa7L4k+PJUnDTB7VxzJt+m1OLLWtmMVS8ASACG7gw2tz2bThRR76b2m4oBLxKNr40uV
wK4DOrZm3dmnlV1aUTCjfFyruUyrLM8+XHxuuEzvdNFCr30LdGXO2+3faRaHUKM0K4FByW6EwdxD
J6TrpQoyRRoDrpO3CKt/tJOR/FslydsbPESwYdoFyYPRjss+7r1VVGOoc1s7hKt2w69GRCRnylzq
ty2cbyTwLmTcvIBQ3eFkjX+D0qIAM3GrBcz00sFF43H+iSVUI0rIprsoN/VchpQw65vUKRyjRCnU
mGF44b01kMdgogM8AwTH5rAxSZeworHTOHHMMCb7jH1/4cCKTz+ABJkBblr81WU4p4gjfTCdqAWd
mURqRpNqlDLtdYN2uOuBp8mhFNvwm9n7k8rkTjM5Iwri9RcsBUZMfz7bOg75BaY+5txVc5xOJVVI
uZPM18pUod8H9Ow497P3SBHvTUnyzNVY51RFQcdkmrKrNfLXjnZAhu6PDLPpkG/XwiBZv5dL7V2o
JJfRdU+C260Lb8feARXA2w2eupKu5kfPXF7j49xb06BFk+4Vuaf8zlrLtDIcKKLfa2msL7qhqFiM
f1xq7/tSe+WFqNnlOcUkfRWn8KN34xpSoaTD7+D6cYBwdybhQUQzg52RoYZVjrFQ0UIPoYiN3GFN
DBr14uZ4DbG/4wIWZuOWNrkFSLuTzryOdodOtZRy9y4V2I9vsZdbeEdB6sFnOt01JwQX+XkYiAj2
zBRZTUUed+Mpgmw/MXGmErrUmEGOi7PneokZ3PXzdF7CY7Q/HrV+o0lWzOH0vf0a1qeqvyth5GQf
7GheX1ovY4LgVuUZz9qIJU0gE7ODjMKNeSuratn/Jt3y5U06LQokHjDuZdyqf78+WnCOsGWtyNdx
Do672Neeke+pThFoMmy1u2GAVknmBQYJmzkwuCuNkrf4HyWe6RZtrgcGiqCCFFlqKtrBJPv8DZir
6xiIAmZw48Djkc5yUNQCZ/cyecz1JN03le8FobQGYPuzIcvufLWIyqgim2E/L1PxnFPNafwZigP5
M3mMunv/9C4EAliX3H9FStzH1YpeADvAS7T2R0Eo3J0qVfj33TB4FkOltHhBQhb/2DFpxpN0OO9w
xdfluHmnGU4pTixyCugTNiWoWOAsFRnpNU5lN85iBJKPKovTTzvWNKDEIVWjalPpbFh9i6dCE0LP
Jn/ithyH7iMSI6LxdrzmJMoVTawLwDJl5n8XMwsFQqmh1HoQ31xxvV+S4aSwqpFZsKnqKXvRgUQ/
Htg/fYw1erwf6Xkxi3fvzVQEkJ8z+5UDlRJ1kjDsLhnsye1z0lR0mjoaRhnjFI3jVvKYYfZVI28r
Q9cBck2NxpdY+gDs04G6LCioG1/hjF8O9Qislwivc8ofWy9u6AUYpPpg+E5DC3o92j4tP/CYdjVo
Kik6Q2Rf1Fmhkc/oYoMoBpKgsroa2CvrORaOo3GUuZaa0N2Tpt/WAzLqgtM3s/gWC5imhbwuUD+H
Pbuc0Z7S9bBGZWBiRMlhb5bm/oHTT8VHkGuPplgjlQIRERCb0/t4501SqjpPqdTAk+i0BXenEYum
Ws2ZgjKMn9TQSpz2KqURYy4i3sK3XSV9qVUeaFyoiL5HsO7rs2sDBla0a1fQruXgnTMmb0nEbW/4
w5AIWaePDxQPnRhKQCJNlyTE6XbuWcIDlVbxJ3K+gXSqIhfDG4s8+Nl0LsUS8eyAi6Imw/I2Srj8
g5R73TYO3oCu12+lYuFsAKj2xsbHAgQ+reXHu/pIjoXrVZIiJD13QIAc+NMBsbuqqpXEPqjF9Axw
oHCCGkOIQkl08RlS9agt9YK4GlF8+Im3Sn2As+9sGd4UwpA5PpI0syTiWSYEdqCHWfWb5o4L2MWx
eEwHspts6HE1NUVvRdEzF5sJu4xIe8vRwpVAzA1M/8K+5XpRg9vibjVaF5V6xaK1MPLujHRrE1sp
lkYFJV7V+JcoggIf0EpCVzghYfwE1ZAVgCtOWOmS2cfIqxLWiXvwPekGZAh6H/4BFFqKXyp49nxQ
E0kkbT/fvuYi8MJBD6nMyu2eky/8zh90t2OMIGA2KZmRGgwb5qzj3fJEzPo3uezj6xk3yXH+yP3E
fM5Wq03ZDfzGq+hIWtwhFniz+9tUnciyl+GpgfbC5A2Codoj8m4iQPyCXDwAmIixhte82mxSFZuJ
l7zRy2SWwNVPM5Uh/E5PZTCkB9reDJ2RdMQK5GkidsjW7DCNPJ1gHHqGKVW+vYkekLgxvtLpB3z1
epMWzw1SefIzm9Wn1xI6QbYRi0NX9GuLpZm22ghmldZuJP09eVmBVuAJsZF3ql4KStbrsI/FMqtQ
RVhoV+zw50V22l4JiGs0blzuUf+37kalH6bqMienA5/WW9TjxlfbWWHyidu0lJr3a1H1Tlc8FGlP
GMkjBIpKurxMw8a04embYas4ATLz6rTURjlPKJcDRMHHfAkkE7zxZC1IGyOE58tq+18Nb8+G1ckm
q40k8D8U53SWl0ZXsG/TyeojG2mxHmX7hJhYMRC4m3uFXsQ/MFAi1PkSTdOeNV3gMjud8z8Y9NBX
XWnz29Mj1NVhHVH45Z3Z78NKzgObY0mAZCDP0jixwnQqdDOIQMelIWmBTTAP5tQe88rK/iBfNZaL
pSRJGWGxSMi18WYABPE9cT25aHa8TjujX4BuUEu0uOe2VIa7lS0QsXIJsFYt0XwGDnMLFWGVVMPd
21zBpsXDJxmWii568VnXHo9kYL8oEN08egyrwqeftACKlJqkKRRVOJQx1sAF4r6moqm/doU9dcTc
mzIKEPyFi8wZoBiGygAYGMHRTzvSvfsIYhb/8pU+rubfiWRJlMI5oUq09ThwLCAngEruqzPcfTa6
TEuJezfOgfYzSRDgRNLraOCbUuV1yg3WMPIPvaGCBSWK/jMyDUfcdn4Lw/6HOVypJIRAucSiZUFK
22GoGn/Hf7k7ugknFRe39x05oA/jg2VshXYf9V6B/GnUM5YP65p0xGF5WdVX7+xXRa+SrB5sKqCz
WDpojtgNVlD1DJpRQqkpPKgIzgH294EFoZ1lfMTv0YGOXTSwNFOGzOssyBZv7tyotTK7iQrZF5hp
bDG5Rk4AW8IKa/F+NH7HYUrJuQl3lrHzyQOaL8cZNKsSFxb0K3f1X4TiOEtIIewfgzWLN+fbdeiD
KEaG7ccS4Bow5U1vH0TW6MuejJTjXbVDg30nIgNElVzpqlzVqs1GRKZ/afaT/nQJYOAEexXZPzU5
1tdki4ryd1OcambSLRZOk4+hqhb4No455QbOmcfDyNXc1Y5yDAGgIj5FCKlYGYLzk189aqm9wt57
RnRehYm27IYl/LNYt/pmhyfuzdJwO4C8/u+5TqtlbMTsF5BUJ+rpIpGPuzkMlovghFMzCKKycgp7
qPM0nZfKSNmQlrpgkcrpEKma+8AfrMqbvIPTbvFOvaQussqNa6Lx+k08pM2TU7Rv3HKgaFUQenNx
/e9J+FIujRTInwPxSiJjE3/rfp74kh4KUtEFcpoZKfXvc3eoUaGQHEcDMMIxftPuCCNQ9J53tKSr
uzwZg9rQAZlscxF4TaI/U0kZNFv42eV5QEjUSatEgNt7SzQer5blmxXjZCdTe5B6EWVjU7avy8NK
VuqZv+9Fnq86ixHkQFTMPjeQFS1YkG3NhNnu1Yndfu8MR///xj4fRzazrbpu1/dnCdHh2KaL2W5B
hR66Dc9PhPqX96+UhlnURVBn6yHoHqSwU+eB2Dgo+1b+EsCWNVc57RBuNFmLBoqoDZ6J7Je2+4jq
sNPdxR7ShyW37ijYphBdzYTlRvydXLJVOrFNejdGoSRnR/uv0vyyBGiHDIsNny2W4YLHqUyDh2Ev
RqKAVrj5/Jk+87lhxgbHmxd+/y65lU+Naitg061d+2Gp8ArpRs9IJoq1C1oN285Vzk5l+gPm87c9
jPVQZ+LXz5E88cJ8TDd9VW/kX7KzTWxIL18bW7RuyFxQcFXHPzkrg70ce6OT9B2AWlMBcYDvMe85
W97gBelhUsBEun9PdeVFO0vx0JwO4huULFkPIuXkJH+AKtKvF/yg5j2i8CWE8w6JL3inKt8Rf7b4
dqC7hiQNmnG30eHi8FSVlceHzFQu3TwTwWNWNQw2YI4jWIWWza9Aw6iu4MhulHxEfgYWnFWj6VIH
8qNhyiIx0uTh/UJtwWGOKHDmY8q1QqCLVSVzkqvoiOKUV8xzR4ZcGl89UMYSSbZUendqJBDOXSYX
cr6V0cbJeBSBfBSMCx2rGO6U8H8ysKjmy4rTuSk5y6ba3uZt9ths+iEtbMykuNbfhJzY7dxTErzw
m+sHmlUx2gP3k+06A6v6IbXiiDCCT1SeDVROuaBZkdwXTNeQ/M7kKeQoLejntoQoa/nDMYUwtEMq
rhevQRAbBv/JbkmIs/v+8yW+SfBabk5Ixf+8+PpLtfflXxqhtCVbyn4qFAbF7DGL02VHIiJelna3
AZS+Z76ganeWMBPD+1aRjDh4jlNuAjbl8TPPo2PZ7rlMKjevzobMhI/wlsAREdpwZeiE2kjutk/F
jpfaGMjotGW+4ng0aAQiOWfYw3KVjQpD9tBr0Q0lSOMtffZWi4x9uiVWzpIpNkcd6nUWDKftFHI7
K9j63zQkV1Pia2HyH0HYzrDH0ZyAx0l9Ud6oOcu7NubOpq0/qL8OJzLlKrYXUUvh+eaBOD238vpC
sPF8Qe+fHbdqDi+X1LQuY1tMA6//FICST2qxWVFUIKK2CfivYWVD0jQ4oDyXJoCcuegYgf9aRIRr
Us3VNI3r8mlo5MRqq0Hd+pOcV1+NXkT1ovpOZG4x4Dz80DQTnxcyMJvBvczqazjdQhqkYJ8Q7i0w
iWhknlrrmI0+gQeAToBHEvBkWXTo5nWtJDUIauc9a/TiDfR44IsPnNGKchP2qJ2HVUTF3eFfxoa+
GPw0veGzw0DId3itTUKNKP/sYGdb4rUzpLLaaFMKnLQesNqRRzqP62r+bpVbnX4iHN/eCVcrWTt1
/lljBaCEtb87ULJ1P35VQTAAuAQ83Ma23VgF79etdGoIuaylEhPsy0Y2HpzNMl+lqHT5iQdnHpK8
r0foU4PtoK7CDmDFbJn3SpwV1iVDXrkVc1lUwCqlM+nYlNkNkQg8ze+/gS+uHzWmlD7+sN6ncHZa
xuA6g25aQsLtlVuGZqqOcTkdCnAoy66Q4QYkDFW+rCG7XOJu1PRouMYWH275+8Q1q6jyFpfS8k6h
xCHBh7x3Wh1aygYZuz9mjqN7E1fHK+x1JoIoLbEYJZrfs/pkkTISgdRQ/5+i7V1BbRc1CTXJ2wUB
F0g+wWoPi3RtpZnpOeUqzmJlcEX4rT9ZgqbXGAQdsu3EywtfQkkwfUUsV4iyPQssiPSyE3nvZUYn
PaQqfF6oqF9XK851sF/alNKF2uL6H7uKrvYSP8eYkxXORtHGmZ7N1BCEwCdU/Yk5GWf5TI4fcSur
F8QtkWyJGJRdRapxhwwDlQ7xf807PmsMvkgUaKWqmrkRuvxKztCsXwxxw1B2jarkAgYp1v2jyiJf
mh+jIcB5TATswF2k7IQLbgvQ9um23bS63FVOhCAkJCnGfQjC3wBMYH+ErnahoXpEFKurqd6qIVC0
i3+bcT4J+tfmENISbNs3OmCMyLC0F1zD8xzKhHmAjyHQjPFgA/DxL2APxbtBwolmEpwk2AjwofPu
/qC81Bok+IIE4QB8qtO63U6BybRRuOxDGLzlyq84mHYDo6E2yCH0l0dY8Aj9ghiHVphZDoXI4+Vj
2cGeSrW709J+eJUOR9/5lih7cBwNX2Bb4AVhCdY9VQFipvxgBzdSFdnCqPJ3oA3E8hhXqS2Kp3XH
ZieB+ulaBtwhKcaj1BFsRWO+8J+uupzmEKezvvNffSoo52E9VbuYfijSLT5QhTT1mLVCPMU76x5J
CP3de+BtLlXJ7T+ZzCYocvrX4J+5izGovYFDbiS7E7i23239NlGnKElBFTQuaXb/lILqtnbViDrp
Db3WTdg/hPpjbu9zyT3rrdNtV3nc/Gc4wRti0B4+udyp22NIyjtgTLFmsd4ohWh6hLiIoCHknfIz
3SCM7jMmZiXocxO0QA+tfYDN/FgUmeLNyoKcOJVJ8CHtGIU2efgfHP4YmkrxSxmzoQ67YmWbV03d
kaamjiGw+jPmx9mpZqyWXVn3LKkh7kt5wDkaNlz2CPeNbDPeR4zIO1p/OpzdvX2WZP8VvrjdrfI2
GsuKmawwycj9oaY/2PtgiRakYKicsIcHdwO8BH670tAvvkpJP2/IhEYiGLNL4tB8kX6+gs4CY0yp
xWwEHiNjIRfHD6HquXnHVqtyAfV8MBrx16ASlMlcX7I+DA8DlVmnq5bmXWwwITBZiyBO900sUMOZ
cZzBh579O51hOFjsjjZAtNKSqCpXqR/6mbf7/oXFMaisPj9gD7Kofbv5vNULxgxaOknsbc8RRChX
cL5VsORgFolpWpU4jDC6yMX+mKExJZCnHgA/8o9hsBqbP/1fQRa6Q6wYtXVZQ+O18hTEE/QB7dvT
MzBBJx0WYEnLvPDmSwpoMGlobgtMw6kJO+Xy2vlBtfGKSmsLw9HULS+JrV1wzPaJnAQ9QyDl4h+o
XkA+boyBr3F7yrlGwtgIqNMVtEmImOk9iqvUoyOPm1hQRh55NYEPtTVsp4MrL5Ivv2RvLXMwQVDW
QzKBDAYMON3fVs/6V4YiTkqyEIRbfNsdqV5GVmev7WjtidBDYVriEe2RJZHsYFHKWSP2oalzUu5v
l4bqaxWQ6bgucB3tA5CxZKxmuFfGW804rrpHgzfScpih/WdZnqrJjPoZh6ueRwfR7rdhXbhOG9K9
FMjmwEf1FjaVhDImrmsRHtNy7H+dvmxNdR8PZvwHJ26bPj87MRvbnlHvAeFVcPSjSoRwXeMcIr0Q
SRKBv/HWahoK8zCeBPHEVxPX/5sDe+56Y59osTn1gQRe/I273LCMqzdmEvM/nCr/lOjVfXGmmUV6
Rh2+nDvJpMxdsnaKg5vW/f8dPbbFfFXzSamhev7qd85kF9k0fWYsski+bAQUzsZO3kcmyHEkBt5w
GCbipbFEE62whz1k5SBJhBBUALWw5GJu2Bx8BYVymm0kh8xfw7fXdHeY3A8GSVvNIrXp/NJa9oei
7ZN5+6Var/Ivmi+JYC7vlWyjLWvz/HIYcqYgJCf6ViqxLB8fIccsghtUo9dogwUaeEMHmYUMF1Tw
TVSpI3Af0wxApyHQ0eFMQyq+mAovy3Rw7VKY+D062063zPMsA31bdGcURW8asG0hhXwXn+oTsvnV
0egmJXrB0FXjExPFNQuvgk8qkImZqCvX7LOIFhkgQqLG3+UfYUfrQILklMUxLX+shHUbAkYvp5Lk
GiPhZqzlRy+Tdb5Al/cYQutVrIWQ16biiLZE4RIgFA9ALFBmtXwPy5hKOdT5jHLhN+uwdgPj7T5x
bJ9ZEf/xuAknaOp2luUtsMkX9nXuTRIDpKCjB4v0AS1X1L8sU8VdR0t8BdJ3UYiU1QtabH1iDlLK
H+ZZ82ekUgJh2uROHw3l6D1DhVylnFnIZyT5lwJhmXn6qc1ckamS3wpxj8ImDRZNYhNni8f2o8hK
S8uuWD6ERGx0e9wqGd0+x7XGEmAs9QInMHxo40fWpOoQoVREF7PcRWbqY1cqmBA0ulZmkhx0EO0Y
itONl2ypEaAt/rOLfwZdZHRglU5BIfABypEWoDKset4MRi+NypRH1Q/NVwOXU0Vf+C0xAHgMWxh9
RCQO8OudD1zwSb6L3oFno05FxrGGUPGtaAuhKchFr5QqKDa73JPVHzWqa35b77t7B5LSiVZC5wRF
/bEMtyjsHB+nvYrgX0h8sNk2OtX11vm1wvU6tn39WPeowwpH7XnFn34mqZj/qnO7SqOZnVyoD0be
wXow2v3x9r9Mg3/JTxb+oZpD8IO9cwtcKPVkCV8tMUk4AKGYacVYW/XJ673bkd8k3NHmhQxbPm2i
s2ZAj1Ujm4TcA9hujIGKQtpMgVYWYSiiOi4hGCiP9lq4YVJGdlxd+2YtNB139GIhU2GBze2rdP/t
iNCzqlVKM6JFYdmbTS6FUR1Mz2HCBQ6mVX2Vys0sGBp1gHS6Sr+6EqKuAWEAJAU0v6ul+7EfIXgj
x2PKfWpBgPZdFNknDvOw5un46ZUfDf71DLVizh9MuxXZ80p+RDgYE6+QTJ9lpvkMBEluTe2Z+4BE
EmzUSYXUPLU/9qyf1MNwWMB0g00zEYQ9FeZYdF6WW4pDdPaVb5IQl6+QC2z0Uz9hTHRjMelJToVU
9egG4Zibb5n5XMZuZsUQMdAKFQdtzN+mLG8trw+dBVuaAsm1QKhp0MsfknoOpmCGMG5g3VQmZDYG
TW5z4haAoCr1kQa5lyC0hiNkKzJ8ZQTk54WAqNfkre+USYSl0oL7E0WZ1WQO2oc9s8+sG4/pK0NW
S2btKWdPftd7+0aq+9PxbUHyg1xoWx3YhcyOmlr6HzQq7WY/zVde01XsGMOTmLpnJm7pxcPZfFPv
LMDGNcyt9yX7zJBZIoK6h3d65AUfp5FY7i7jNfz8mWnGdsIeHfc+oW2ZR3kJLjmPIGbHgTP03FD8
ULawIrvD77o2kMKtQMEpVMBogEP8M3IlBjbo8HQlMaOFb7pfyPeaO4OEfeDVvnrsJT4hxbG1e6w4
7WdR1ANo/7wJcJqdAd75GzeOd4OFsrCkuRLaQyugdRnDOhrpvhK5+N9AmOx7A58T8zkZ2ldURsAq
+V0lnCxilHG1/0AGmiuetQOxGVqTK+G5P18gwsqKzgbD/tFhnntLAzTFql+HhIj2O4oA0fSjeCyt
aZrCsVm3X/qoVZzVnWWlFkIcMwj9BRJZhrx1W3P5EDnVmjG/955ax8wPmbmP1FFBP7t9D6T1BzX8
JVwj2rafHon0sj4veLXH3BnSvytmvzwngLUMF4oNFYnOhxrHWzxAAmmZb6eyuroCpJMzesxUoW1u
twQOSGmDvqZ5xsq7YYmal4WhkWIazLPFQRLgMAk9Iq9n2ujRF2aPmujoqK88QCXN6Rt5qE/fbdXu
sd5SwuEvgv76ZxdWb4Fvkqy0wLpUCJjZ1WB1u5QuPnMiWbFCm8p7mSLIVBbVZbIIvA5SUIWu8gCD
ie5JRqzpkyTJlDULt5ZVsjfNTcQAn3w/MUScn5/RiXjCsYTzlSMuI1thm2PUSTqZ8N1xmIvkF4Zb
yWPTx/KgySyFFlpokMnDEg4DTg6ZApVgM6xSYf1BgxfuM3y7m+wf+thUDUotnCq4ckzzHpKtteZt
lo1DafMq3x9Wltm7cMTAJRFHAAaL8Nu7oR1U/UBr6HqwXCwsXNe8glWBHt4K7u3Cal5Gpe5jPbg1
VTJv+m6C9IgfIMZvHW9t4LI81NU71N1RafJFbKqvC58/sDh3zh3fEiIBe6qVCAhYmtjesLX82tUK
Hd1qoIrF+PBGkQB5INCZyTaHLuRrZHmNxb/7sNF/ApLUBugu6+U2UaALNn5/hcbkfQ+1ihH4bsI3
gRL9v7ZUzh7wZube0nycklATcOWSVCJtiLawq/gZMOTEveDQn5C5zYjelujjlhmC4u/Bz2JXSfAq
cNPZgJqWXDbzpmjz2abVhoit2N2t5tpnUNx1zNVA0UHqrzG7AB9aBxsscuooGnYdbn/cfL24h0cr
bTjyjLAcIk9yWBhXDXA6xJWruHK6aOCrNkCQfcyloCx6QoeMpwNCkCLmcn8z9JBQw6YeHMMw8XiO
R1vMjEpk8yjGTxFrYSLda90FDmElsnbPB8Gecy8arkbDdNolaPxAeL0oP6hpG8sk8UKGizJj9YTx
3suEJkAl5/7Y/dIzRi4a+l+05+lTDVwWOcEd35ZN5rQHP0jFKmKzrnl4A0yx6jSRBjwfYYRP0EHW
e1ybEG8rBAe7fMkoLsAqY7fkRcJTzzBungL7IRcg9samCWBZUOpaQlI0NydsrkqyMISPayrdyQfQ
RmrtqOUXxpZsz4LqrhSEKOkg049OPStaiDYpLMsBb/Scet46eeXOKpfENrgvbPU6gE+injfinSPw
saw6BVik126wQq/h36tQhXemRg/f0fo6HaK4ZeMmlJSADjPwmZSZYrqE0yl9TtMAa+Tp5dERdduu
TocCy57P0EmrojkQgR/VAEWH/+ZPbHSAq1fv6/jCSlq2/W+o2yiG+6iMn8g8XuGzScGVNYqbU9rZ
UXO+y3ZMmSZxzB+T/NxsF/zFpFXnVUApnfnav/ripTvXap5C7huCxhvA+OeVNGvihwbIz5o4okqJ
z1irAIZbwqx26z1IcUycVWpSYcy6mR/pxf2b9vzx+ETxh5Pno6A1htwCYmie8OF5FyFQzyk8REDt
JbcCVBre0Jb0aWO+G9rrBd3PpX07mxQwYZQ9UoBXA5tj0wWHrm54tP1gMo424tOsB/aF1SQXD9K0
Q4R6Q8vAcQUCnGUgK145MtMRlYjQfbZFGbgJGVdEE8bamDnU3CujLfSC5ljSTGj0ACbYbt1ju3Tf
sKJwLWLzoVovslSxZRVBf7crxm9pM25RCoVnZIZ2pwN73faM7ipQeopX6aLmf8lZOSBDi6EGsOps
leN4uY4PF9FF/OZ9pH5j951VGVbJkOovmRJj9AVKa912MSHJwqWR7k0GKTbhQ7Ibn8ZP8yzhmJL+
LQ4VDfOXXpYQe8Hrt5dvOIVH2YG076xNWCdtcsNNy/gSaBtH4cjzhBNTW2Qez2YtsxZBYpee0Gik
W98a2DkxO+vFRHERANoxE4WVpZSHA52AS5PN1ygXtu2ZbDciZa3n/eHedvZktkdo4hZ/gwTu/7yY
l8FAJ06D3WQiJrXe370WcGnJdnM8muGIH2g7f9qxf5dwJ/lzguWZa5w4FU/IvIequosut5odfJy4
1tfvHuLUZHY8H/US06KgPyz2DgOt95nlguG3FC9VqRNiIPDOJoeyln2kZECfk+jDqz3CFuhzVdE+
ZckX3zFJ95SV8/if3xV3ZbSaz+xviU7z8oTOkkgC613ko62V2jEvoGhWfWncLQHJ71+W8vR+MgKr
ZLWBgukt4bZCs/U83e8W4z1CVLGbdkG8XQ3uTCKLrdbhdlQRdk7lKXyQen6teewMwnaET0R6Iv8B
hR7bko+QUuIdLxvXW1mXHslnpqbCb6Bq7x1nGZxP+WnsumKoJiQMk+aPPDE+p8JadEryseTaVJp9
9pmIbXMVkITA6jlK9pFUJtt/qyArtDHciYz3EqOyuKlESzXqhU/co75Lr7aawc6TYxKSSsl64mzP
UXRS5Ygrl12+A2QJW/NORyhn8kzVUHMBIhLq0Xi70gr4dnmYM0Hj0UuLJZaMIbbZekWyPI1VeQQk
nzbelagGgPthqgXEgRrsagEg8qilQnKObzLHhegfCKdRfGCAAVPuBF+cj7p41wvF37AQs1ylR6be
dYe8zrH+CIaudpo9mkcdu0Rm8/Id08BaAPMX4PbnZ0rX+S4TEc+oIDmrf9Cxjxhme4bEHPWNtB9P
IjCjtfKrsUHq8kSxh7cC/LufmoElCIfwBp8+7CzLOX2CuW1zlgIQlxCttp1KUc8ygn1Tzy+P8rFc
laAAQXokTn8NqBHg/toXcwd8RXlRdlBbkHvTGJyltT3yuVq92+cKr4FTt6l+Z1urXjRLd1JuSvOJ
vDPhh7vN8wBp9McqQyouj224zY6m75k1w2r9EFFvScdXpltniZgJltxxlT5OcwAT61fEoNmkx71M
6mDHBBwDBiTiuqtGZIwOuyQllwAEE3pcbZCMf2kBdIIqAldc4tvFghTy9ge+ymQq9t0hkrhUUjEx
U7LncU319EO/FwHzRksFmzCg/Tn/wzDDvR/X/yDv/yeEcueHM2as6ry/XntMRn9J39q0U4NAoPMj
bsYMmjjvllLICLsUSm5XUFFe9rwelPfziJwuGofjuK6rOscUqB1op1NB0Kj6rCmSrcsXLc264NZQ
0cu41xqQCYYQSwTlUfVkKHiqAmVfGaNSj0OtBrLz0q8fPRo9q3A4yYuma4uKYp0phoHDt8lL4xz7
l1T01mgj79LinrS970etDo2+Gl6DEsc9t3TXDSohtHN1wtYkTGoZnKGh7otusZZg5a7IiJEScUSk
L1RTld8BJMhlC5Dgr//IBv8Mjl2USQb2ED/5i6gJiywxvAuGTKj2sn2TGPkGxeVHv7iIrD1AbcOb
eOAFr/4w/HxKYj4iAIfSVRZ31XM825QXOJFxQUyjgw/kRPM183Br6rNxBRua72ZTc+iPx0bCxR9y
mEMOVadErzMtv1fl3C+YEczAa7aKTUY3FxGzdf2/miEMssyZE99W9pHSmzV8oDNJ/yZDd2fxEW+M
oOicssCeo1lZbR+SZBCk2B0bIu4/Hnnbe8vxoKkIVENvfW/E8VzOKnJO1HGrAr0guYKDvUEVWho4
91QeWCyzkoD9PZg7tsyF/4z06AmN0B+v26R0AbStt3taHtlf0GbzSntCeuYnQO5gqhQgmbDie0rP
LFflELiaptifDkL8iZ1WqTr8PbbFeis9SnT+1EziOOsPcfa2ELb7LbvZbStFhJ7FIZhlL7cTRawF
9lcnruMQE5AKAFlJxpmgCuwqwjdkJRNrtByfk2hwTp8JAnCt4FtcQbgnFT1eVB4RiLiPjSashh4z
cSfOYW3gHWiTGti0Fo4+RjQLcPKKurDa4W4GemZ00ndE5UlN0BVkWFGVKjLNgNf3V+vB/Yhp1YsT
a01zHSdv2eN4KBDQwvvsx5i/FUUzyDiKFsKEKot/8dZOdrz0aTlaMiP8Unx+YYkW1gq2JcRgI6qX
ib0p9Y6Q0kIUfB9VfE4lffjKF3DR6Pk7TRGM/RZyNuQQY5EMkNatp0bS1mnAh1pW9LwLhaMGOAbg
ifCscOmyu8B9gtbqgg34Oy++XeZAKtYkD4RCJtKPpWCh6ZTb5wJ3mvY1tbBCSQ9T7qkZsaHUVOjZ
dObhhEVD/u/Ez1RBMkC1dLYbr+DqyVeMfYv3tH1WDa89vvv5A/zmFqOoRP2RnzPz6q7j9Cv5H7VC
G27Oi/5sTvtcQh0tSwfEUW7ilOwp2Mh3ei3S2Im4ApfHpVBgVK1TiDMlws3ejcBVo/j40d3id6Op
RPn3wN/znv3T7FThqAWjxEujEbCkUwN0jZk+GwSC6/ah0AG7WzvKiy+Tkj7r1E/ZYzc/jDq3ULDk
sM7TGht4E3aUaFDrNWOFDbM74OHkdbf4wJliDgbBe0qQy2D3unG46l9s1NVsfYcAveg3P1/0L00E
VKQ7DQ+B+Ycz59zBK/1PKMXJ9wwLfqojIPkMqkbb/CPegKoZURHooBlRCsXNuAkFNCh1n+t2YjIL
2ibRQ4FayzqmdzFcY+wEQVDX01iI+fEiBmB4VA5Ru8eYawHEY4cQW5JT0JX3V4P9PUNtTDTwW9qg
uAWTn25WP/gZVhknczuN9qPxMmy8SfD9Y/oyl1kr0/dW4j2yuArmF69SifzmsNTTwhAVQBM9oBJj
cXrK/OFa7h46JDk8GhHGDhnfqmpeha9brBL19rPf5OJLk6cx6aQEOqxEpa2Gwig0TF8rZe02ZozE
ii0mYy+3s51gBU1EkcPBi25TjfIwUI2wsmpsBpmQyNdR6ZeLrRAMyru8MUFSIvbM7bRzSYQTFXsn
MB+9JXIeAx57k+jQuN9bzoCKgyIp0N1hE43GN1sENTCI0xxc9ZiaMcH9imudD1RQOSGjwkN5rVOT
JlGthrFY0RU19Boi1eFeJlClgK9d4+k9dK3PAVASkXM5dfiaJVdvq3UrXheAGDNxSCkSE96pCR68
eQetsh8twOec50ISmAfEGmNNtu+B2Iork5D9vOgSUy6VaL/ugyBu5DtInpC8YAF2T5eFUvyIqLkn
Q+8XfEaCacmUdb2Bfgl9Gqg/qWwfzpvkCc8Rr8DKwPk3Ozdx/AeMQTDdR/6w5TQbl4Zp4FoxxXtb
/+4fTr/K/X9ggEhFgyNez/eP1TTtvHm0YcApJt/+YDJomJ0k4Kq7an8koqH+4+5Hsx+6uxlezQEn
5ObBsrKPcOhmowuYHM2I7qAVTthQx+7m7VPDmWD5FlPsMNW/X/ffFwGBEcXXCeZiqDj6Fikgq/lx
PgGIO4BUkDW5D2e8NqMth6QxVwwBZzGW1PWTZmJPX5aKWwoe1DXCzvMKsvwZKbjI4Jd1ArzK4c/Q
uOTM9akusjYC2LiQAgop5tKxXOZeofwtLnUP/J/KoUGhIEKAsbV64s9L+dXVJYM5C4ZqJIXfvErT
di/+eGA37F5YlQEbg2qshE9s6RfcXD2D+UE7/oI0ggv8z/NKduznoxUtMMm+usDYOPgngpUN74gQ
yqFGsJgXHsQoLy2Jjku8zdL0bq9gBUyEBoOwKp+Xmknbq4hv856zA2JmwxOM/kYnbwEFLDGmwLqo
UUim8xT537YraAqydTClpb1WrdjYP1a8zOD/rd7yehq/U4HD9rIE9T2XcKRGEfW0PApSt/3MCfFF
53lEg4uFxf2JZHF5bVJ0d5LPXlecMInR0ZYrek7lPH3+cP2605aKGqSXV15By5/Q0O8LVe5Qyzxd
Hq29Rfrq5pBjq7z9v7fMTozSzKOWy8TbLNwzSN69aRpHwCNz/7HL2jj7w/muIYJIoR3fNfnzW8sU
ofOatmbMies/llwKKVYz4e2PSQTCkUInnfDc1AuupF1sPQZQvWJ44f1UV6Kc9pvV2nNdJv/dfSUA
3WpqMO8+UePzOGRcW+Eii3yOUQWpDpaagLViXDLE+DGxNLt62+Mj9rfhFCqpinVJrBmkJIIW1DRK
6ayJ06WXLONyoFO2mMKC1lt4Vv86AGP8NfMmSnhlQwK6wbftAzPiU/Fv91YkuwEIswZ11yRbBbsk
9HWjlecLaZgtS8A60+G0x0tNw9cgsWxYcknwQeLaX8aQiAbBm/EarfciW6mxW9Xxl48b4mX7PtLM
2Zr1Tck+ctERXlzlK0uXNsXpACiCOOQhpQIREVU6ovk3rlk0h9dIgFpsTcxyJilHOnBLc+I1khmp
QSRqrKxQNmNqKMf4V3judM/Muqa9yRcDSIZrhG0X0WJ1KSVrW9UPA0NP/GifUCYI9UseuVTajaH9
cD1RS9p42wAuNrZ2KjEBkpU+tPMmtbRp2mvoOXWLG7EF6OTcp9ZMeDqMT7pRBftZiOBNTa8YCLzl
2ngiQ1r7j5eoqs+CES4qxurgyOzRuZJkXbyzJw2WkVe6mUPzEXPRLfdjW/1tCsGbpgU6jxwKFMHa
E7bHYZ+5Q+vL/dtnVP2Z8PF9pNvxPTtQWgX9DteNJGrLYCHCRZ1Y4W1FCXbtDMO3h38uSlFzUO3E
vPKx4+M6aPbXzJrVxdZ1jmNQN5ekOiU4wR6grHb/joareTfm3ldOQDmJbjbG9ghq3032ud8SbaGU
ST3jfzPKFcAIPnLBWxbDux3SRiGuVYYTvMwdVDXOlYxxkReUg1S5dLwR0dF8rLBrV80DRnD8XGNI
1vSo5/UTXighfhDqB2NNmAli2CeesH1n5QYiDh2KMxwbHNjTkO2HzVH7lHb00px7w7lYye1keizM
i0j1shMGai6MOBi9ONFNnBOUCWw4fLy/AYO0ALaoZ51sU43UpIMaImqPfg7imkpNms1NUN5wqIpu
ilNjtXBy8TvB6uq3CNAQlfjhKyzw5kht99h5BLmQkObr8gtJke3IpFRA4N6seluVTBCVSp96ndmH
hzJjfKKrU5JjZ6dnKJVfhKXNH0K4Oq//7UR5MHTYFAKMQE9XJ9yaeW4efnsWsZ93/wQAS0/7yS/m
Q7Z2HkAlsTRaONfSkqvAKnzlk93ntPHu8Z2JMvKmqnaIBGZAEKi18ntH5eZQpYRb+l0iPXEj1A5k
MgD09at4EYW/6HbGpYu+Ns12sT5f6GnYVRPbE0JfwWRVsp+6l9s+0RpIyBXufAD+lxa3c6sTyADm
haF1r48+OHqqWLbgaX2OktoHRBuZGwN5dMQP1Rufht2rQebjnrMVPCVzm8tuC00G3e6Fs2Rc/GIN
lpKh/nf29uppNfO9nYREC1KArr3KqDkXWcCYBuFcYIPMVMwqsoPxvSbIBrmr8CyjsW4WvITbtapD
3rO5Km2DT0mGOo1Ye6RjR+6aqvVu1039QFFy4k4SWMO4NAW4ySEufkUD9rCG5xMF4U1osF68VhOr
pe3nayUnjA13DKHlfQ5maQ5jlBYwO6M91yMa8TyjS/icQG7JfYNU6305WHyBA90ALNxDYfzs5XJb
484kvoef/sMI2a6SXN9x2xXYsmCtgs2k9FIpGd5CM8C3KnBaxOggp6fdpalvg8vr7DSfiY/a/GrY
1etr/id3Fi2nhZqgjQU8nMX3N3K2Eanw7CFHsVD2+JGSrnpQtM42DTRjB17bQhREIdKXa264YI5I
6U9/jaeh7CVYfdNornqS2IpPQhJ2Z2z2kOLyrFbRiO+sahYqv/ANW/QpxxdNhJh8CEo0Sh9hN3KO
4JqJfTFeYyxKrMq1e974dGmkvQX1CUo9RTgFHj2WxdJuD9xSiGhMcjQQEL5jksDNm0JRNRtww+k5
31zcakd1YkNNZqUuEyoTOHLMZ6KKcsK84ytU14yj3HE5wwzKNjhvMSI/GeccX3RDbAxYFusGMXLZ
RBsRqracV4JpYXTvyFssq5HX0efYn29RkPY4G37z+TWKDo0Kko+33QioSShSQ7mV+tYgY1KIxpWG
awdx09v94f6NhszZlUpEx3vcUjtOW9Mrqt2PrCNgohfo6MgRGazaWh4/hEzlF4ib3uwXLqHZgsSr
4vwqKn1/iH7FLjl/iFnl50b3hWUhNsFt5q4bgyvoW1lmvtyNq/LyAWs99Hw6qMz8Jl+aBI3rv7ZP
uZ3i3vs7M50Pa5TPO639TM8eFihnm82SnmFGprCDS/wB92QwheKLTrELfvse2PVDDuw1hz5ZIM8K
Aip3wtFk6fs08+4IPDIeEg/BcrKA2b+QNv75X9A/GPSr+itDmM+XX3AI5YtMp67b18R4xQU/zSJB
R4FiIek5M0pG/vMN8x099hG0l3XrbLKUx7J0dxqC2z5OM1oW5c76GncOX1XlvhteOfK08rMfImw4
nLnH2bCCZH9gEJ3e0Mx6jJIQB+MIYAzZ8VIclXEHwaE16Qnzq9aZJwZE6z+HNnWLartZaaaZvKEU
l5WMITt5J49rQwKLuSttmjGIkPEi4XpuovrWLmaowEXgV71MATorzoYBXPzQIewkUj31EoKyOrJL
+iU0aPguvffWfP5OFwXhIU6yBbf6l6TcI81HuEWc6b7TSxZyDV4ELRkvOwBhnMFyDUp8XdLwS+DM
B//k7PhQz3diua3ICCkt9WthYzlN1RVv3/Tj70Hq4urEQtyYPoPw7w8CscsWz22qBuXsw6LBU5T9
QFmkcYX4WTzwSe9QqT3qgWZNIX0NT06rSgsKey/H3jwSYsknpNksjevAQMpROsm/Z9OGD+D0HE9k
gMtXFwpkqitaoo3vtlVuXORDiOqGXYTXtQEYEfgE/NXmyAvPqkB90UyNBmP/Y/nJHtv7fkSEv/p7
UCxCXYBwzEirTloXXjX7SumqO++DyKFTFzE0Krz+lshJA5evcstrcHgvvyX5e6v09AljGkVAYn8A
agId9FVxtaGmMi5VAk/lo/IZOsGxIpkmawuyuv0cphYHCAHjuZxyIx7v3EiiMLEFN/FvS0wvP5Sq
Gsta8I17nv2KYUHj7LqDLGRbuEuE0uND/eKnalr2ccR9ab6tLMKmn8qL1TNGPO9/z0skBQwigJ1r
8/MXahds7z7pFISpmAZCIlSJbMWXsQDh2Juj9nuDiyny4klNVVrGGj5LO7G7xHxV1RoMrVg4iPcJ
+kmIXZVdBjvqoxghXBK2BdNy7DPuoHkQogHqkoR1wbcTlw9qP+/8NlVtHk8e4cpgaU77OurBrDEV
f5mmQQhIvyWAGYyUrFiL9FuQK61yfZ1+uTDEUWvp2yHaQUGdwit9Td22PbULjpO8uGs36mtzgVRH
2E56uXFMIRcZt6lnJ1J7FKcDXtk42RDA8iAmqKQu9etUAn1cBvM/kA4ND+QN4IUNiT354xrYWry8
ABS1eRdBExztBenAvOT+bhGlVH7GgkwMHi2qxKr+W7/SfCes/iq3AxuIlSh17WKZwAthm1CvGqe2
tyMLXfSDV1CxDcLdXtMfLeBZ9UDLPq+7Vq2KXPJYE5urciHzYtCys0eCaCQrw5TzWHcbFvDSm+eX
u0xGNgR2hKzDYG+v/6o1JhkDvosJ/1Ft36W1EFZy9jDZsdbjzjxDxosi3TXlGSSEmiSNV4RY9nSF
a2ZMxS/b/+d4JyboLqnr/VTmcf73s9FmOeksxMmy9yoQuG533iLpbvkKy8GwmpivdlQQ/RyX63D/
jJUBJYi+mZs7nwJDOkU6q0fGMzS5CZuDBAn4aXegUZvWKuGnBUXc1bOmg742WSJat7owDIu9ZcKa
4ZLjImKGjDmp6BX/g1tdn5IINnBfUVCQN6I9agayFmRspLfv334x0RWnc+3EQGEPrm0CV/Py4g4e
JAZtVOVBMA3JXLlXLznQvCbqq40Jl/RaTJToO4kVEZv5H1scqZijOQnAGqreBRQ9Fp1L8p5rTCsv
mkGg5713cEFlkWuDN/H0cEWv83sxvYyegKzrTCCL9UvxJmS1ayM13sSCICymYOQQ9pBVbKozm7vf
NGdfq9rp6IkXxayjxpzweoneWswqI6wcr1AiaevQpNUnSEY4mWH2LGEhEYqyryznIho+tbNcTifp
Q4GhnEBP2aGexWFTHKtp6S7uzbf4p07cFLQvKUnOtPSbnucozxw0S3Dp6+AQcfmnRha6s13nZvF6
Ra5OINMuPOJJsVufkBAEcIAgu9ADlDjBSBTmNyAoemc4DpGgmoriRUGr3gTEdVa6wtOmYul5XVKT
scDWutNGsr4pVXEBZa0KYeBorrIQczKoXB0ct4RpQ6ybYZ8zlJ0uzsQQR84UlCvcGaqEdRG3tB8g
SZE/qj47YlDY8FpEwp4BXC0k0OYSmZnbbPujMojFB0wkUwObsJYp3mHNG3nUGVj719ZXiSzW9gFv
xIu5Hmfz8Na0jzf9/ZataWJoaSv4qRkD1/pJEw4gMYsKIDe4bVNe/jmRLwWx9636vJiGQmAzCLuL
C18PZ3CfQuW+GNaxz7NjyMD6xi8BnNUeRQM9Y0ouv5CuUXNaLKUEhRr5rtfQm5smXmR+DYFMHQM6
MaexOIWR+00ijBmTKhrR0ibxLvapl+xoa6jJmsNCEYU+f/dW8lodYjcsBw/Yif3qDdoD2DxaTvyO
x8/r1EtpAz9Ksyqbamt8DJaOfrdLnAu7IiBYmDb2oAT5CRZEXWNCfQkM8AMZUevzvOIkbXyZZ2Yu
GlEStsqgUpGHG8fN4oxXYQBz+YZ7goUMm+QdcER8Y3YndOTgeGJxFDZ/My+RnC12ilx1GkABo2wi
yRuhBzjqcB2U7rcvd26mygNSWEe4+JEYVOxqep2edXHheoqpc9vWh2ukQp7SVsZil4MSyiHfBryp
09cwdwYdr6T0zFnnJxuVY0zO5MncMIcPLCNs6IOVYd7LrLPx3hwtBXh0XkvgbhFXVXZqqFCPK6HY
UxsQJ6B+G6Msii4WhePHvziZOHPBctlu6nOIHkFkvKcbr03lXqbCqpoMVVklIsts8GXXckJCkLGH
SnH5bgkMpo6DcigV8OfxzicPSnktIjZQmBrY7EtmAJOme6uc4zfG0e+Mi9t/PgVTUskNkLyxk12G
C53wpLJEcopcRgMK1seZMeesMqWmyoYiAzHPYZu1LdeQA1nk+Dg88NWfmuycnbFUQJkDnNa6Eldy
f3xl6m7Yce3tHPpCM6ZRS0jD6NAFCPnj+l4HODiQ1m/ZVd6B0J29sh5NJpeBAN2TmQ72CL064Mqy
LYc0dfSMyCp9hSYSpzRBfrpeGC6prhYHuUlSadGDVvNXyx3utbXsq++cH1v1f73nezYaWhNabby2
ctihE3Vvij6DBP49VEYtZTNpd6LlGXDhmQp9txiZ+N1TTD6bKibHPpyvRp9CT9fEq2PKFxKxl5tc
oqr+xPjPdVRymaSi0ZXomNK8mcOaH81tDxTutvhytQRVAHjS985vF51+qyVcLTbajCMcjE+VXeW5
Ew88UJdPtXAz054OO/26bo6ujz9bTVMoX0rklOBnbZAohdgfhVOF0TYuGM5PxMwbAJ+0KCqxb2vP
JNixlKxzCqNHxMdSGyX72NbURTebOSzjlb77Fv4YIerUkmhcdChwA0XhM4nM9SuTL/Oo4BdrEjhZ
jCO8ACjKllVPJQkBjiIrWCyTK7sTPbNObkqQZDzSvN/MHVJBv0XinYLXhUoDXne6YVuPYUzrulSg
Bdo9nrvY/jCNC/9UXHsKHCBtk+OQ5/N+DGGzQNUqs3NdjSbHgeLIr6P2D2wwcmDt9cu0bnTBtp0T
qeXsBSQTeQKVtg/1GdyFjzcxqopLmr/emiY9UuvNu2psYXkeu3ezfV+6pOnrLIxv78tEuy3zhIRk
lxywOd+20eq7q36aGxuZyQRKpFa6znn5us1eQNQE5cLyUPzkvCnJAnr5fL5FVLkr7DawpP076DBE
7l296/ZteRnd/pAf4KvAjufrfvLcl0f3FCu8v0YS0H02JC8grL6V2vUl/86MCfqeG90Ly9i50Y/r
tMdUIPIf3vSJtshRGmCALClh7/YfxwzQJx5MN5EC3bHWZiLr10kSaXPjG0OTUHUfpGwYQRgsXVma
osBJ+rcu1H309ZSsd2Wr4pR/eAlugOY7NH15xG4WxAPsgFpahrWWEQiUPo0TdicV9uws+5Mr58lT
DvqozBKRmGB+/IFOfKw754HFG54hU5wGSyG0ZB5xZoVL7iPgGZRyxOcHwnNPphV16ZrtK9Ffy3M9
zO52M+cBxBwxCxoHZlchzLBrrQ/V6sacr6lHn+Zr8blLh789Uh9Lcnsj6IVqm2uJ1ZVOp7KakcOr
GkV4y63TE0IyboIimaNgGzj3w6Yw1C/wra38YyLIgdowkG0qXqUW2kya4Cqetge9QGh6GRHpNMAB
hqjIPNKoYkvnFyhe/rLuNe9urFxoJMiYGezKizNZeMioKkGXPz3FzauB3WnmldqX8pcHUHot5vfK
05kjBaqE7ggnQaqqG3rlgZRgVbP+t/8rIFdovyR6brTiVe+C7Jl+jy9nChn0pD+DNm5qygl2guIV
9AwjRPk3ku1llfYQ8E4IeblWJK5S/9MyhXA5CY6ZDTxbftHAOX2BHToPRnXWe4gD8uLa6+Ok0wQa
dtXuYICuz//1mt5tlnt735ogUm7+hE8lv9r1lJe55aNtcGa38ZJFsy1lPgZJhUuA80QoQTX2pwHE
NFgw6cFdeOpLhui0MOgj/UrjrS4d4D6yoHBdCPgNkqBVolimN4ui84QEL/miXbzj3ik4LSPDrjLi
R/WV5EbrFuTsohmAI55eVZXg/oMgy9PMs+7m9RWaJB4yqdCnlPHBvd6j58Z1zvg9SS47cTp1MoRO
dTNxwloDr+EbY5+mE0rsKQDxwgG4g68mcb21OJiHyrq5dYNlMijvIxfsWPwLMig74xauZwkKlwq8
Sx8Qo9kceFTYvWTD3EX6VJwVdSfgcr1DWfXFtkCi4judKNIUJAogqpTlnbIpSrzzOru2DrZhmhMd
ODCTemSIp4lCpIAp4wiEujtQd9MR72zNIynqjkwMLQGLlgTDA8JXPKUWFcRQXprbMWbiwoS/Lztd
1EniXcnqgVxssdY9jtmU4HvIRYtYwQTKtMimUcMVFEt/0KrnMTZQ66Za2rY1Z2IMfnauwtuydVD6
8UHGWGrrGBzwlfqdBcbnGNxFE65mMZdLYhAOHdWcmQl41fugQmJWK/pYXdRUJVJoY4K86ThaPOSF
cOF/PPegjEcxTKm365QNMSjalt7BoeEV1vzXWPWnkic4EDVdmC3yWhcPXf06q0aASR/DYzFWJHpm
mHhkuulUNrwKn61u0RTmoMmhuv+y5cJPfZTJ0X/ilUeROTwmKavlIe/f4uPHma/VkemFDWVzvcNs
j9h8cRiLSK0L+V8hNoBY+hR+oToHnEb1TYeS9mr2i6ASnVd2CnQJUhfxsewG1YB9k61dNmNMC80l
OakX9zOVgu/qjUWH4J3yjEyyj1/ial17gsPRo4qJrPP5VOgMiPyIzZOZc7x+pddnFlSTIwkn//PJ
I1bltN8bGkDnFmt064QAMCX5Vpc6ecjzwYoxzsZ3kdR5kc3Mp+a6Sl30L0wVfTvW50dRsdrTbchZ
svNeWVRW9iMw1OsioSNdvjveO3W5UBVcM1uPjtsYPNofZaohPdJz2WN47931WF0Z7yiOwKGhFyCB
XX0bd/qaUFwDF9Vq+Y06h3qqGgM7JSh5ROm88oKZal27aFDesWum3H52HjoCCOm9pzdww7rnydmj
hYKYZqAbm2Ow2BqK2hTuroCiA7SiD9oczj/wfX0DXVoWC+PKgH6YuLzA8BRExWFzzJpi25NmQZSl
H1WacgzrXW40IRlcUGQ5Q75LCoEL5+K3Ql8nN25eCfTqkABo71ol71GRMsjiZgEJwhVbIeaeU05i
ON8InepdnSlJne3hiijzWDms+gTpvdE/f3PBgtoT4XsHwOxcAvS/eX+Zm8Q3QuaFQJ7YM2C2iiHU
NW6pDlWs9Zrn6bMLpHhqEut1XKBUYt3MqGALxpKctkqxCLQsZ63tOq16dTHvrljw/dRNPOXu5ATR
TwrvvHhnLEOUrA/l7fEhPSzcPf23xpeO1RdzUpvRHG1iWKWa6c61iGTvXlZ8kj8EymScc7gh5jL3
XHaOAQJilvt7QqY55TYDxiPpR9k6iRmRg9u6vExuPo5NJYhcsg7MxfnIp3KeMD0JrjnwTJstbb8x
C8ABzPzMVcxIbk1fVgQFnWTxawxp4JyvJwKVnS6NuKy2HD3tcQfQpPx7EjzEeQo27IrbyqeUCZ1l
mquvUJoX5Wkv9A4EtyDh3H9XVrjwsvQ4n7yUQaO0oKF85ZGrebiCOj16/6LijbzmBMziRHUaZyGf
WMOFpbUPMMO5DkmAmK/s3mQxBICtqDaKzxa5GwCbZ+TMUdoTb6RUkMexNdYJqnVjaxu1YlPv+RLH
brqWRhQn8GcavcA6fttoEK0GI5cQJgbbXz65pesRs6qKimO0W/bhp5dtxVBkcUnHfl34YV0iVUmB
IHq6BnUCay7WMFueT+c+IzZE1oEnp2siZqIq3X4ktAzpNN333hg5Tw4VKHYNQKkiYW+GA03v2+mE
b3aNG4qAE3p+8je7sqfntO1ZJHyFsR2AIJglsLxs67/SXSOl/SVSAGGKmkY0OJl/RVw8WYTRzrEX
hdGuvxl+il8kNYyiBFTB1APKe52VwdNrNgSLdBoKGX7jaeOsd90NRDiACJpGEn6E2FvfPzRE0Ano
aRvv86LqVWLJFd2N3Izl+tPkuTslNUrcoUYsR21tveegzXZ8lP1z7qtz+F23QEc5zcZv5P3yOIHy
+fE7BVlUn6jrVVvk+XYOXCHLzdRx9MCnhMiakMjyybs4GIQq8713AMlfq/KpxVEg4eJ3de5cJiFo
yrrdEdh+ub+hTa1HgU6ApAbS3T8ATEuA+36txqw5HpuASUUzFVWvdkErqBvqkeSzeyyf6EloftDa
dAkfR+XX95xtXcC8SQTOGEhLkqv+uFdJD0pnNiA/HfmhE3EAXYDnnUo0clQgfidWzDXrWI1NutAX
zZPOQszQQRAo11oV2jbJ0uU1tZd2kL/GefP1Ztd0HWBCzvZG0PVoyIyiQFeVeb6BFesWZUUB+tjG
o85xz1XT/CoD87ts9ume7ROeC0k8cDqpjNOnSOgyjGeOreUegz+g0XoBt1w1GwKDDOrq7qjiYCsm
9APvpHFfJbnak0fe97C8W70Kv9iP8TgjVnwQJbpOzDukXufQnjioUe0BsqfoPL1avkyTLjiaFS2o
GAZgDyIaMyqjLHYdhPgo1alWyCJ+WkkWgjufk1ynoyiVeZW5aVDYfb+n2sVNdde8HltcyXwYjH8V
7TvmyK3F6Ae3ZATcGKXwaUuoa8zUrikJsDGXzlYmvn1G3Ne6FCl3RR0/Cz/3yoTKOvItcbZpBPC9
GewX8SdGUTbGP+22T2wU38tC3Zezq8V5BosCAlMnSyi5iwPmaN/Dbm1RovqIYDtWQj5G9mYkOevz
h7jgQZGHhnh1aQEVkNblTjFNW4n9FDLmvY5ByGlobeoslFhCmwEaOLYQrYFT2/lt7HM6OC6JxiV/
ZjdXr8afiLIGtUA5d2Eb08lDwLKI4dVlNVUez8/lASshEdoioNsswK32nH2zQ1riV9EfmX4t8gSE
K4hlYlJ36ngq9DWaEyrQP1QvVCQA9+s50lFLOm9eCeY4z9hKxPA965OnyzHbtRGgcOf20+EMaEBN
rgSG8qP6eXzMh/UuxgPC18uvmoGR27TLS6BlAf4wSD3W+MV9GaMa/RiE5CrReyHDtdMB/UzNdPNI
OftGM1SLL40CNQNyzfv2VqRDov3EJ9HbXJXl3kF1BgeQ+adpfUaL0lSkkg3l5zbRqzwBzBwaDpTw
rcIH/IvK0pQNmlUbnBL7YWqiHueKplNTNrp+mMcbPCE2iI5LnBx4VeOY7B+lxNg5GibpoJzNIBHM
XIuPcLT+k7f/zccOAwtPk30JbUUgYyiIyDMiWzqzpob7gtzwzdXQZsYmOSPpYayv1DlirK0j7GB5
3Xc0V/vgFCa4TKMgAuGljfMpQaKHwREl4UGs/8fHabiBXOkaXttEZmfrf/819VrLGRQWK/xp1kL+
hwaua00DZdgY56maG3cPmS70ZK4XSez6PTYckk018b0G991/lVTqox9bPZOmecn8pzlSUWBbA9FV
bZ8+hj9Gl3fgSvxH9X9YsK+A+xeD+vI1bDcBt5lOBeNjxsyPDpZI58e0xDNPdyL7CrKZ501b5p4E
I6UiJQrEptrvPk3xrPN7sMS1Esj9XJIGDI1x+sBIPdYzI8d8TQOT3s91yyJfYxxJ5RPHgukrFxnF
pXbN4+JlUYRT/xsKFEDGy0h43mRqRMXU2WP4phnkkJJQ7uXY/WHjFcgQUiatxOikQAxOOY2ehTV5
9oLyJYHd+KXyeXcUwulfgNgSrhkwbSAGPdxrMM1XIsX2n0Z1SxcNZ1aKAHWCMgHRtgVEM7SSC5Hj
0WMVpla4faeWjYNUyA8YvM7FSkPQJha07lMDgPEX5catOEBbdDoQe7pn0X2z87MUCcvnmSRerldO
oB2/tGWAvAR8JDINwiA8uFPLdFlFuq066GHYzIgU4tATXfqaWDcNAjzWXKt4J+Fbs/1R2+ThSp1H
S9C8guINAsHZstTftFErIqvDUyxRjtu4UXaywmWNeBKjwJiNYWCDlsa78iddxZwPH4KWN6xGct/v
TrDbv86Pz30pUC+r0JYxj9+GIxk4uHGqJUcf2qdWqDuC5eY9Hoki84HbSHAEVTBVKMvzVXLAMspl
03cTe4ll93fg+YmMIKoMXtndohFYiMg4SgYLfbWRS0h9/mi8hi2TorsOiZD8aUiD4A7NWvE7D0Wr
GUN5LPUIVSDRZo51BNyKgmw7BCzJg/3IM1JgrSHJiwHq5YReoBPS0EW6St/VzGhd/12/add5qdju
SCOw7XY7aELM2THXQg0ZexwyRb3dDJ/fE3a7hR82oBXw8Obp3VROW3OWJ4/18gbrU1JcF9a4rMtd
7zWzmEWTvLRr2aCOJ3AP3C9mW/w5HefIc8V49PWD1WwC1Vc70FhuLHFE1FXyRllLCJoXVSPcOf32
q6aIenVPFRGn1++otFvoCpap49KNjqIafhh22/P1yd77PCfdBkAfySWZO4uxuZJ+kiluoKuuLJBw
nuqdikIJVUXcwkLsuvO0H/+w9HUUpOVN1n145bnY4qo0fA5l9W803QF5maWW8qaUkmplblLJ5szQ
T8eO3qN8WgqzzA1bLwsI9zQOH2jmtSPlKuQnwZ1tthdidxUSKHsG2gLHPHYFf5bBkSZIfHjYzV6n
yItY/oqHkX+vQqZY/9FaC315ff+ZXAC0cE4oZbt74xocCdXZjzlTPnYdkDIFzozjNHn0W1kgBRI7
DBlWm6O8EPW803gqQ4JMI06BtvEGBLwpHP5NWkxpN2PZnNKKpZikxJNluxrdi4rGBZjlSXoDfkvu
F9FtbNG1tYWqX6w9ck4B4BSE2OzUc29rRTa+d6HNymZQDwoFlB/P0s5aYVtZiHkfBQPmzvZ6XtSI
1yA5Ri6ilpK/9/T+BLo5RTytSwZ7DeS6MmM++zpssqI/aOsmGxPnPaFA5muS3ajfj+0b6LBR6QBt
h//rYdmbRUgK5g/sqA9Tf6m7NZ4ar77GMXpZgievWx2J3SGSd6kgbSHlSSc7un0GPsWdsFg8NOSL
8n+Z/zPsREm+9EWNmIMeCRJoZmL4NHDoA0fCPvkT6PfSOmM+BWruosQhFM14n0mGGWv7xgZIyTcs
0fFfHqREv5JRBk737qc+vLhIBv0CUsZB07flIId85SCrYjIe5eCnEmGIADgJcuLa6us1osRr4YeZ
TymR+5Lpme1F5Rz1hm1mR7tk79mihycZ2sxBpj4ebOBhe8FMG7xZtQADtLIXCuxZOkFZPyPIiU53
dXfQuktDrToy94HcZSsl+qFtpe6bRLZl8DBfpstaxdHBH2uF5uArs8GZkzuAa9mNhuaFYql22MdB
jSp8P1uMsKl1MQMIqvBLEu+dE9HYz6vLihV7LdalntOb7vFy6OGz0an0hY93cVFz21NSMXYc+z7W
SI8ZavPdtI33Z/TxZ8fRqtvhyWfkSZ3ZdUirFpbAvxOfV5Cms3CXo4tHhwL4VJPa9b5yHodMyfBq
YdyZHO93ZRcCA7D9HAR61q58UOrlOLu/91BnH2rccrQ1y7astD4hLH0T+eJS/dFQlQsUU5y4MZrW
sKdT5k2xDoNRgpT1dQMEjdI0/uThzik8TWwZhfh7zneHtsQ+wCEBKb/mQMmgM7KTgAEeseQTp4Hf
6KsD8XBd9Fhaa9xp5n1EXLcAt62c+N8pqzpuHQo5Q77MXP1M5485EEUr6chRjY4PEq43qV/WUgBo
DXiHm19jTnhJJOJvBo491poioIa2HAPatqQd4ClBhVBmghZ60ySYotR3b+oCxLFcP0w1Xox7kjsA
Crh9DuHeuLEHYOz3uz6haaVmN4pgcBrrNehfhW257ppUt/Lh25J3/PgQtWlf/2EKc9i1SK7K77LX
Xf4YX8gHDfddi19G+wycNIAgdFFppQ6kLCiEV9Kidq5c/JajOwiiOJI5PUg8ivhghRJ0n9n3Lww/
w7ai16YIoZbGGivhadz4h8emCwLwSLlpC6vlJOrgUUjiojzLFYLgSFlzGCeUaaXQuFbZLEZ23v9z
g8ZYFaZBcTnCHSYDxsQq4+hieAcg8uyFmLsunNLqeHFwzOzZsDJBz8kayhWkd/ZV5fK9I84xWUzR
neR2erCMb6Wigdq+6B7yksqW5vTX5mplj4UnW1HuIOneDfV2NHFmOeELptq5Wt3MbP78jB0CEekv
vQKPgdpE7q2njt1TJP0fFikCYBMgC17ZtUW3t6ab6eplt7cf+squ58QjXvkQiYDDdYI2RrX/b0pT
5nhML9MP/gdehTTQq6Hvi4nGzb4qb4C1Y1XBJQw5+peqatK6oBy92jvERky2G4y5O0HhgI9nl1sX
yipsXmg5ilS4ngbglOOcKWgaoU5D3WO7077GybBAi1nQEcAWWosuFrTnzySlpzlBXBjxPlOg4fRt
luqG2jDo/GqMm0eRa9ncYwsxYknxuHRZVpCZo5Gn0K+kZYbDkDtLb4EF9nrf5UZUPB3xXkXWH4Mo
AJBCYcFNNfDjwdTNmPKyUrc048w6brF7Qhqv/+wv3CTsAWza8tuOqSIsNIBNCz7qe+9HSuWW98IC
04OhLTqzpevDKggk+jbO0v50pLPKaX3nw4UecrNUNs1ZBhClYDtNnBkSFVfzMIQAoXsHVQCu1/E5
+xUUjBJAA4YOp+8VjK8UEMUXPXn93rZYR0gmDWLlR/roYcDpfO655wecSPc5unlt6Vy9OmdO39CF
WPqMnI/mQmifxqoqkn9nWPWRp+xJgpi/dKOohLsAyhz3JJnYSzDjdNrT8OTvqATVXlO+ZuwY8+gX
L3ZazTf/FAjZ5xNXsGP5WxDNTu712wF4+pOm1oi4T24E43qJVenaME2TFSXV/7PE1SgwX/Yz6onS
2PmdcV1aFTi62UquDemn8XlZeWO1ENmuKNAEjJ99N0XhwMBmXFgu9Y4LNOx+8dXba3Bp85NALAEb
8+t91MJ32jAyOsJ9NsZ731yz6CQ1rk/Vw6C2cjSVFnU9J0b7Os4m2hdTmcZs8L7cFmBka2MUHIg0
P5vliPirq2U/CAPVIo90vRGVwdl5141/4PP6KyU8aMClTUBrRIjGzxnt63fdEsQaf1kW9kdbZ+/W
nNL4copdJekxudc5yIm0kXJ+oIHwHBynNOQFIoztV3rqxbPNbufw7vKZDdzZj6nKtKKLnefUcM7V
S1WmaDdy33viw4UVpq3KvUHOuV3nsRFxUTLQJ5fmYvN/+/I4qPMDyYzuuGJsd/F1pyAda4SnOtnC
GLGZNaWoqYIa/qgeVAmWcKXWk9/4p3uIZ3zmLgpEWkV99N+5P7T2wschApfL+w9nWDDqLsL29z/m
cWHC4frhV1dfLVTHixxHp8KzK0Zc+Spyfr+6OZVpXrVZwubql0Lw0tV9PVdb5OuU2ylts9E6qpLe
P87+w8ViYxuefUXl2ntbI47qFa3Zz8v2EC5Zuyv9IqAPtifhrnqn+L5zrg1bDBclGHEJEF8DJhAC
CIDUWvtpFyvtuK4QmdKO7+YlYcIKvcXK5vFpi4K2SeGfPMCXGarxjbwcyjf9TN2SVfGlg8yFmds2
QPsCRhi+GnJGtQwwKPN/iV7mW0zy2alvRnpkksa5gmnprWPJEdL1ADis+5ZtzIaG9y6n+egmdotp
j2EdAJA6dDHKl7JmflIHO3lgP3/A1D7v5T410D152WsTLJCxwU/p0h3sF1Vw63hb4lgFWGRSc6EU
9byemt1FaryeZVz+XkBh/mb+4JgV1NozJfqgqssLb7B0RmiQbytJg4NmIkscFOR6VSIs7i1bYCUh
6mb0a0nd7GL0CITBzCVdd7GOnEJ5vWbVjFT0EioqdyIgP35hlgNXaA+l4awqsxnUntW2VKYW9o8E
5zuKfMYgFNiSb9sRCPpJ+v1Nbfa9xP6+/5EPpZPkUlLstfToNdBDYILKEgUKXhni/v2qW+gAhA3p
HfmA9KfgRim426QY9sbmCJmoXAQ5tI8mQszCA+ac//VVv1qKj0tKsAk/lQ5SZtqO198zglU3H+EO
3L35zvdSut6dd/zrNVe1Pcvk/fg501xMaFA/eJ1/KMrn/+9syxYg6GpOPHbmdUP9qJFyGqYWNf78
T0Cgctym/Vjrwb5paLAmIoIW/3O5vfBW24cQ4roSPmcHllKLAdJCP8S+3IKXRImRgZkolTa5NJVT
gn5Ncjf5MsNm20yb1T7igAcfYRaIuG+suZGp7crOP7ajxz7vU+doEkD+3JChJFQNsYAieB2eK7P5
HM9qQgexOMldgyqeEE2UJ984NHgdGultwTDWQA6WrZ0gnGS+0LoY/arJonJgVFH+PR6O1Tv59tcm
jUrEw8p9xg3POSh62AmafpE7AyrKre1bQlmn0xtWsOcZrW20Kt6Kaze56LmtPv0rtjkK2gn4fjJM
+yZipYMnWKdhx9+JyogqKONZlLBHA5k5NcKlmLWyU0OAsmr9AWdxZ8iu8haes4hBvS5l/CQeBDek
cfaTK+u+CnATAmwKwIH1LcF03m9mOn54sVmqGYU3DIgJOA+gwbjEUQHFYTpGMUcdNBbN4kghEDrJ
343FbNuJWqxAfuH2SS4ms6qX2DinQJmLvvurpihe1FSnqA6lVAISVpOvboLiE+RfH+HczPMGeFJ4
16mBSAhXTCeEJP+FI0Y7R2mrChiRYTSW9v9BFZGfXiNsfQx77kkySsTYSiFZTum/a3r/OGgePazQ
ebfj1WVT+/pkXbxkviSWhcSqAW3c/+R0KKtcbpJt9Uv60xORhqxUdzXt8p0FZBt/0KuQmigv0Nkl
GFBIaLXGJKloyix34xLEakG5f+FjaegCs0D7VUgnbQsCpBYdishemS6cRBBc37xA8uiILL5ZZGVr
TW7aLskavnYGJ0sdYuqQ6yKKUj7xzIxEKC0ObkLVlF3CSnJadbQYxbo9OGt5yxFwqbUbK0EJtfQa
f+q0dRIotO/1J21MJlFQkozHamZhiBCQrmqq5FLIOZfdakECfgspRt8TL9nFEvOW9yDVcdsVg0d4
Fxm0ct6D6p2IAsOQjtv4AUd9ePo1p+p8dqD2en5lpPDL/Z9P1mH/NkOXuq1AQjnyqGGnKQjska5V
qEiF3tRt0mtma+mxtx6bQr8MDRy1vfST5Eq218ZHHoaDjxpfnhWjutCoD4zj+QnG8PRZoSPaHb+T
aadRHOjBabZQXaWbufBefh2WvXgcB4hh4HuSM8vWmoOkgJ/1gnPp7xOrALCYOcjHS4AmM8NZrj+V
qWf8h5rke1CjxOb2oXnXDNAijDK1G9GeqPL3Yu2N2DDi3nmUcNeFtJ1mppEFRMauVRkgMkBVUKus
PDrt8y1rYVxsTJ3qFoitEqf/4El8IDomjzwu8kkX7Tv23r++1ji2fKyCKXIAuKWyNcnTFRTMT7KM
AXU2eq8qieS+DC+GMbGdxP/jlo4wZGl7JScUquNUlkbnCyz327hdXSDeUmVzazMlvOKtd57eoGpH
x2un4PCYvVqixaV0ZAEMkGc5ZqLnobS/MNHPrAreXqLBYpnRZMh1YOWHjyTRz+akR4E8BCSycGYa
5/DcREnCDVwN/y3Cu+JvpOInLRhdAD4a1Z32PxjTLVaNY8QeSyepfjbZfW0nCdoYaJXVUz4eiae5
xfQm7IBuytD0dAIlnBVoz/tg/PtLo+7D3fJFGzay8571F8cQnj5YijUREuZ19NIvF9RbLVhPN5n3
gxUCWU+L4e+Vcps7nW053vlupcK64F9aB+CXKNaDCQUADsXeoTCwJwOA3YOMcM99ndPaHIdp3atU
KAs4S/FCVaYrA98EfC2nGO7EcGF5YwbFohcCpZO1XmVuOQjzC2Da3bn1WUTrx6j382G24OGtlSHe
CJI2lECt0lDDRA1YnnIyDVPPEXLT8rWoZy4w9UmPk7Ev8abIvmvfS08Ghldt7Ni4XPGSN51O6a0M
32bWvH8I9kv1fUDEo6Ksev6YannuuKiyH94enxZ5+hAKqguHLbTz7U0dMICToT8aNQNssbJMTG0K
19B2bnbkukjqGBuemJBMYffhe5iswltbPYo0+q2QqCIG8GhjWaxJwdTPmn1KWIBROauSMx1QO9Oj
E71YvEamwA7ovEe6HkBNmvCH4/xSsSFXH3vLoJ/Ly1useQUqO68t4rko3Fq4lyduikwUj+jphae6
KteaSvsmfphjNzxK+ok5nnpeI8fNuR+PHM1vxL61cSgkGpxaseXNJcwcVvc8svj34onK1jR6/c0t
Cc8dFTozIjvjOubeGFc29q1Ew1SF9u2hgG/BjNy5sYs5X7qkMicJCpdwBxKL+Qlm3zENf25z29Xv
GfU105eIlhW3TPVbR90Q4szvppX8fhcJWmsgfwFYofJ8rdOXcGrCHmdDTigjDGytZcM7n0pKxNa+
ns89rauLTo+nqflZSQKt8f03n0XD9A2ZZeVET0I9APr3ewuUY0Ob/P7CHDxEQxbzlA4kwWJp3BLa
K1DTY942/MEQk3FalNaO/r5wHjf/Zw63O9jmNBP86G7ntEZfWw4bZ6DJD9hMjdLxyvZYAHy/Mtjz
Qdgko15FH8bDSQueqEhh2cunKPDh7Jl8Tdv9biviyOe/UK9+taRvQs6emASYMcjIe3LDtq30mnyl
fm/19wJHZ9RmwSUtfy3cKqbGJxXO00wpUshM/C2gjyTFLJQvmQPrcz5i/JQVGKSGQmNPVJhrfabC
dNOtBiYWlHNtgXla3iXmdhCTJNue/RtCj8RR03zBWc5zuBCYM1dmWdpjLs0WHiMuJQ+LgX7i7Q3q
4mv5iHCLza+q2oj0wmycAjcwL177qRDO1Ox5WtWsIguqq4s6avxD9L+YJJzawxOjqD7K4MkMHOgc
ZDAuszggc/AR9QCoZWhMhfJiBkGDnBl4pU+9lQT7azLOoOOiDgJ4hJIgmj6tn3Dth/cbmZ3jYqE1
8z9RyVYIb4qHatkYKQlC5Tm4qqm+N854yMDlJeyN2Mqkx/jSDvp6kBO/c7A3d/usMk6PpBSrFlNR
IOsfqAgdaSJ5HvMlMGHSgpYMFfBdlgEoW3xRdI1N/Tf2U2QesdTpRUopU0o94iVPiku7scYH8Exf
s6hQ/YIM8dPpqQ1SkvjE33E3xgwG4Jl8lORL0m/QmTc8HOiVar5JG2zyHdvNDdNhdt4toocRJ1ZT
YjnRZuqqwrZ9J5wRKJFKdugMvc2boSCzkDWORNE7uivMV7wlPh5iLdUCWMkdpf8e+hzwki0wLsJF
RuqY8cBjOMHxUXNsutyaVhqYo4+/RqWaOFSTnR8CW1qHdqzfV59krXnE1pxXncy39uj650MiaEOX
c7OdovnQ5Blu9c5Yd8A2MbwZup9fYuSKnEGkZLQm+/SMmL8nG3id0LUzzjT1CFwS9dgMzVnvjcK1
gXspKxb1LN76Atz77YjqefrQUTFIcm58iH1lzlEbGqciCZwa4mArToAF36tCYCta4xGzkVrUy/zN
CVxGOeh5Rg4pzoOlzrwQ2lafaFsuKZreErexx6qk+K4NSXdIAZ/P4UNe8utyMvHfEE7aHeIeji0/
9XF66WnlIq7acvQ/LcyBsffyAXBbMNmdAeBZkdhIXEbeIvpwcMAVYvAuTDftGL332yYwzFMHuLE1
uPb6B8yaOKXfeVv1TnV/OEtRbRcwvVo4Qmym5YpEQsi2x9g0gpkXkjjKXW/70AgmPZzwZbifyhpa
IXFT8Bz3+SspwliZ/SyaiqtBUDmNdi9q2WGhlEOD8eDfXAOd3IJvtezkkOelE/u2f8ObWhxdoSgj
EFL1+2s7KFIy/fHpQesoWrdpa7G7mumeLzIAHPFix5yUg9mvvWkZNqvQvm/XyLsMMfwMGiokmkVq
zxgIWSFMWFp/SpBGwD6fa1LRDQOU2obspQM85h1Pi+cH5w3irLGz+6k8KBySCzQsYBMldLZYKTy3
MFL/bzCLTvMO2j6oC1q6uE/fKIl/zB7qnSiSNY0nSwX88DsTyt9S96qF6bt6iFxDXicXbmM3RHW+
jK/MIIRiNa4iLoGGTJMdUL8Nx/Xsequsn3wRUDyKHkD7ciUEf8sRw0nWYGnxa6khPrHgjLlymSDr
ktcX43Jg3v/W2HuAJDPvKkEZIeZOlvGcfhebF2iPw+sih4HpcSyMB7VaH0+i9ngVITByitbOIs7v
AW7162kCuV+oUgGs92gY4mdFf24jogII6EW+V+Rwx0D+xhFUA5UqrOF5czWVOiraN00+hh3Ib+Hc
Ukjiflm/dT05991RaaJsgJrEg54RZ3CA3VMJ4d7z27YVks2/6IXjH7J7hR/1u3CDXXHpmSo2Chd8
Q+K00AUbET7P5cx7FQDONSbo5B/mxc5c7R3iBM6XZGGdqlNsFrJ6H47SfbqPJHt7S6h5Br6lCO6p
k5N+OlBA+toIXySYjH/hr8PU9xTftfiZP7xoe0o+3rkOEqRPgRLG639+cSNeFtwY4BcLuX87/CGy
H7nBHXj6sOLbULmq4GvHXAJiZoZERA8pgNp8OuvmEyRgUqLuzugu55VzQ5NvIHMTpoWhJDlelKZy
2LonubrJtckQAmcylycjJafmY03PNjRtLyIrk0CD/QyQ1JtXeUCrt6wY5P4eI4qEU8eXUnHA6CJ9
swGWRTR6M4IVwN2OZRbY3HzglFR/ZL7pKtL2ozRpZBo6QdwnKVuj68hgpLBGkuf+2W4cRDpe2Gmy
vdtF+AsiSPZMBFk6IyShWLqiR3gfqcxju4Bt6JEhvmf1R/u+9mq0X69EkMAA7rNPU2LEe5t6w9UC
6pGx1gJ/tlOpujMWrVyDXjQEvlqmDnfxm5imQT5RfoyrSkUN2TG6vLVV4cnrD3XF2IYPn5omtfQh
KvZpA+wzB1+NzM90q2QFNGDXIoHbDW7+HMOGNP/pAlzQulmdTwKNgNN8j5fqLN8uAwdHKLALr2ZT
//ahyfKdHEbfQJoWoRh6DUPLGqrV9VSHJKrsrlrPP/DsXNOdRCZxggokIqKA7o/PlZG2J7U7a9BV
pgS5qgJYXx/wdg3vaPAPo5AT5Sm8eSrrHAanRZe+VpqVZIUy9WJ2PXQAucz2zoMjB5+Z8Dlh/gnK
VBk9e1MYQMPgDmJ+bHTW5L0SO817OgjOjLnwrMxImCz1AUSkpoSW+0HEwIHm5OWc10IwHrwmgD04
jPhrI2/vNWmZW62KFphycMqqlTZk3GpSfZZe8+fb8tfb91q+bmaNkSZY7con4XuBlbCms8k5uxMQ
ICj+jmDcqQD4zRk2Jc87+mSYu6UN9iy/44avaK7XVep+w1qYyX2wd+FXe/UhvhiD/sVlnvD1wjs0
ujurCCo2ZG+pEdJ6tafb/TcvCkKCypVwS0hXwl0JWIbQt9lHwl4NAzW7+HSCQzqroaVTWDRb8NMa
yWyBZ8ItsxlER/h1+Qb8/hfBcl9pvRkraRYuBdiWFx6RRqt5qqfGuNWB1SyilBfX0lwiVOKGTsTt
r//yuqUAxFNla7uH96DXsgg/ZlS1qO6pQZa8Pci/Nc3xsAeBTYEf2X5rHY5yI7/4cuo7hpESKRg2
YEtFT+HVtcOQTNgKYTEELjU9Kw7HGsNBtug3C27NAg2Qpz7ZLdfmCwNRKo+KLEdxBuIKo82VxuAL
Iw+/q2a2fWTFUvvsKMqPhT+rKHJEvwrW8n6noNlPCNzMjlcjkyN5vkv1Pc3rKJdwBCRbKoxHnMsF
eg+vpbx6JqUkByVmA3IsrAdz+h6GM9PRPHjfGtPQMcZBKvgbDNRNIdBmB5nOk4ajCPPoaRSMzVV0
HUi1NXNwnPz4m6yFgoQlx6c/VxnZHy5iVX74d94nLtTvOjtz8KRBNt6ngScNCBJ1rmS9c7KhMCNz
US/3O2RNb4cKIJ7jlbSknmY/rScT3Riss81bPMLYHj2iyv+PTWAjbres8umjMWU9Gi3OtGPwmuvN
p3hyVjCY87TS8rErjYWYnBnqi2Yuu/9YDaMsH5mp46/jbaw3c+DKaMuulaM1n/0FOrfjazcpKf+o
OCvX+ZFPTDrDXmlxl0tY87W8w+s61VbIi1t05bupXjj2Qzb5qW4sdZE7EvhJ9UtiyPxVA6RJ700M
KFPAhr0d2U5jg7jBwNiNuyT+Ty8+HzAQDV+g2o8OV4/iMjtIHiN2xfEPEsF8E9HWwl4x4D1oEfVp
0ZP51O8LArBn0tNsMSQ/RLoKUAOYU1VjTWUoxZb9Vuf8q0rV73VgSzPaSMgadSNJU8E2d/PxGhjN
+vcqAjft4WdTlLPq+hn/N7ebjUZzG4E6VQj8656uiRXSEFgx9ryKfn0i5RDTuCzfOC2tveLbXg+u
u2rC3bdK6njy/AbwZJCDZFi7A+jZD7WGY2H0BetPf6sNBfKyWcDcXcgbCRgURDBaJulSvt2djTEa
Yxna0z+hD+zznFmAmpf18Oi2mBHUjIXiia9iHPPgI5Id4XSpYmdKRZkD+8LnOayo2wfwk4xIaQbu
okNQJdgVVPeErjwIfoUT43wQ/WwJxfwgf3TFMioMTol7jVMKJTpyAQRHmyohr8IiY6s0MLy4bisu
hjZWoiWBVFidw+ft21qrKww6lQ0rAcFADawH1zHtqbJgxSp+BOFmA/zoMI/ouVUnT6XZAWPQ3TjQ
kafJHoCDoSXRG/Y5iKk6lhb6t/7t+oKpIwSxokZMHFFpv13schMNGVAMzkQQzaQD0bpQaP49jTEW
dPg9FtLvlY5DXb0Tzrt8NxGbhddSN+j0x6LHYBGqXYc8KcxDq7c3OEA3y4WwE1ljD8/76d0zsWdy
y9g1q7Y0vI4zDJp3C5KHjsHHBDlGL7PPxNCtsChcnPDgywmjs8gUbZTalzZQ0RYv8MPkCsTUPSj2
BX+yHDC0HMVhoT8JFYbQp8dqVKZgnw8oC8gDf99aWwCMUhHI7FArIe3r/NysB1F+5hqCLUnjfjxm
gCNWe/4XIXWsX/5DtvVDeCjletI7fXDyHP9O32+83J7LwcMdms+AMHBRTMHu4VJRZ17eEjbFVtGH
kStzzbmOwnRKbSmuj1U1VZCiGbKNQidW+L+UKop3jk0yhNom8TwbmxVohaYaZm5X9E4a+VKv+QB7
4fEJpC/euHJMTdJ63G7HuB0PPeOaK6Yz0SmGVizqHcfAoGXgVaoSanuqQm4Q7YUJ4OJEpMh4UnLF
K4a74ze9MVYDQ/6Qo6VseyK12iBAlV2CtSCnFDAb75lxJy/LZ7JvWtDvU+wh+NT4ZBhhL95Gbtzi
fYZGajP4BX0GodsZBSUfAEgx3ct8Hxlx2qFQPRLYIKKU+syOErGJyhl18886bDbX+FTQFw62uE76
zE31xGZKcV0gk1GunK42UiGO+pvmusiqmmNjKcjT07/QNvTrbjhhwV6x5UEP9ZEaZnNobO5saKPJ
pAi8Zu5dGeoaFIPLjmShQU2ePPpV0H18ntPr23yoPR9BKSKlUe9vJSg/Rvwez7CXdPCn/7tGR4Sn
2j8cCGvOfr7+WXN5m0RhUS/vOyt8W55jVhgJZpXkcTSb8VYNXNrtOz48EHDe2b662E+9VCXALbwv
mk3+ikIW3FESyV5kF0oV20uLJNI5PmOpwDYVqJcCi4mGShLEO5BL2mltpZOPlIEtBE0zt01suf7e
o5kFCRm24agLo4N75GbCswvdtaWMRoM+/4dA73/sXlMI1CyuKW9nLAVqnW/pJ2xsRg5XGLRp+fQK
42v3T5A82ZDSl+5s8C5/hO/3AQMtSc458FuHRXaIJsikgFrLt36TdjwcbOrPVaszXIcG+wJberb6
aYjpLxxwxaYk/uvSUcCIWi0X/noBIUpYvCyxDvn72Lq8QtmYmUch4T8gq4tEUDg5rpKVSmtaeDqN
9vb4wAd8hlSumBHR/YJmBDfAMT1mgj9I167ODRgTJ2K9efEhqBMDo5uNpARjG8YBFjCROavNOz1o
Pf2F5ZTZpW7J0ICEh/UPJmNxKtguX33YYLYDBbkvZmoKcGIY7n0qp8LlrGmJi51QIkdf6WpgQIaU
AHUk67qqGtfrEGkjjiobsGzfkDCbFVRe7Khgd8bY8QGoAxot5ZF2/Vt65bW59cqwLRDPWLqNzMhR
5lMMVoj5PrQTDcH6p3QIh6NLdsc38A/rnVTjmbIlbtlFGVc/iU7C0mDqteoDD7WAsWTtO8Iw9SSi
Ri/WKwg79lFLr6EEJEyc7SJvcN8XioMChFXlx+4jTUMAX0GbZEru3xRNUJLyyryJS+hp5eZexuC+
JNbsssdu4nQ03YbB3wLfrs3nuPK60USzTOQbwrMm6anlDiIFtaKNGlyZTfEi5tNpvCuANr3DZEhN
wD0K+nV1ikE8HOs/bCWgbmZFmdfDW+W1rsCnuvmpHWgDSlnQK9l/xcoPX/9W7GtJs1xu4xgcqIB3
EE2p5EJax7FboF90NXSunMmCGJu6iNZBY3KMZavH9/6qePiolpoMJQPeqQxUWRGs4eiYtmGptRDU
0hsyy9w3N27h62LGwQuh0PNK6Ba+XFHPwFfcY2LEVVvvb5KClk3XsyVa3BBZrQiUu+tK8lyPJwhF
sj94j84hubFtJkcJGNHDB98uKS9h3tSTvgA+oL3R1TlMdIeS9hpsYtUV+BHGproNfO6yhhlx2xHI
s0gUTP6PF+CMR0CqJVILvzuc+0G4LO+U9nI+w5IHh80qHMNv0Nl/+mu3CWf91LYfnI36dSPQMY0B
kCUzXxva4LiKdxl5LiSORHHMQnmg7zrOhudAUJ+xkjHHqsnQm3lOIdbIeIE6p00LN79I/ne8FEYu
gV48MKxbojHF+Z/h717O2nf49cegE5ALRB9h/15ts+gFLWH1x5enKG2vvkNfM9YiG8xytrmBhUeY
Top/rCeZmSJaGvOps3pNVYBSywvFWxWtueuCuaSgcYH1XKX72lsCyuq/u8qRdQrevhSPqIqTysN+
r3k8yOCpSYY7x3uKvNoxUZSxt35d+u+lsk0za2okxQaYA6+XzVPs/whS++vZaoFtLymaL25mT1G9
m8Kmys63RrZT921RsQJOpSBNMLxecDjLbKi1yTk2eY9c5vwBO5e6IRoWXdZ0I2FDgYvXBdJQTS9W
2K8A6S6gcPQfCbjuqZNybFmbtbXpEvOUk3RNv091DCgg2p22L95OirG/pqoL5Gs/SUt3u46gmXZl
xeOo+jFK2l7j4XYZEpRSsiHKOG5S9SBLcKGF/DCt+VdAb8+zbHq+6mz14qCS0jJzWxGcopft0S2R
aCL9rclQsl3N85jb4kimiG8cDTH0je4PYM9tGRO4AYtP8VYhwUohtiEtyTGWxEHd6PamTmyw4xhg
TLXxqvgpfBi5ckgJgDkW+aVcj1O54tD2LQFzselqNbMHI+9oqRuMWmkxrwiyZs3Z5i3o9zkNUj7M
m4sDLJW8I0SkT6RM+bNP/IpPzPEOxm71vefvnt8hfWK/gFNxjJA4ytRcNMA6NENPGjyGOhPdzg+N
hCnloaOennGe3WcEzHP8AeOvc3SRUNjPzjF/UHj/Zt446D5/7blZlSPMupJBdqOqIE8xpysh693g
P240LzISvu4fc3cfIIaquLNCal22SRAu1TipWkLUd9my+s5hhUBgo3BlzuvmXv8dpkzb2ff2x6rC
4BeD4k5dRF7/tBaYz+2uZiTgRFsZr8Q8BIeMkb9mxFUSFfbP5d9jz50QMPR9W3ZD2xKCB3ecOhKW
QpRrEIsHnZwobO76sQx7saRg38cyLjzG6AbDKNOODpGzZcj0W0wYKWMJGEKiSEQ0RPzVd9/b4q6O
P+EWRJVrHQvshtiN59u68v6rmUbC8BNFNoLKw9a5UOClEricdrgASRJhVGtB5zQJA/iPK0ySV4c9
uVtMP2gyLpAai/OeXQ4CFL/th/sDhpHiYAK4DFHEVOqxccPMzWSxBTKdt9xVw8kls0cKiZpOZzs2
SQaXgWSOzbOmpgX0RzFsCjje3TARQe7pCuWLI63FOALEx4KEf1a6H4dRoVZ3td91Wof4CxKrxPdj
zDGAJLEoGhy3OJi12xlf21hIH42H/4oqnb21d7jdgp0wrOiEIUPJPo9ZcuiQHoeLZMY9Nz9KVuTw
rvph8Q29bg0++6Ehu+x5CJaDJ2iYMFM8GSU78fvHGfUp+owAPYNXnK8XJ/G3wQtwVTcbDwENVxhf
VuNYK4Pybr1RglJNknWFYz8hkWonb71BMuHeJB2toz8ukThni0jesO+hBCp7BMLH/MaV8lJmUsHP
PUfpEZw/izKj7zjLZJ1dWkIEVxy+TOSzYa4LMss8DtrIOfCTnWbGBR3QxXftjBO98Ku2jLo0xG7C
8JkH8E2TunAbT/2vOMfKPmSEgNh/Exzd29bLFhIIPBZIIP99OkyzQjCg+G3Lh+kedQVXExkognvO
0SK5HIIQdkeFG4NJxiuKSBibjSOkEcjn2PazGMFqiwT/p252TB2jOQYluWd5srJ8o6C7TLVCOV5W
t683DU1foKRljr2ljM4D9x6WBeTn4/ex1kgI1+AfnOc/3wyDbY2AL9fQkQ2pluHbAUf+FKPsJGbX
RLwmWHoJioQli/KLggcjhwna5QZQkUCLHnrvWP8qbcltm9/ZDHz20yntblmEtEQ27W6Be1oa4LHA
jFJLxC76nK57pnRaVcLitLB3CJQyg+CjjvlYpZ4UIx0LOOsy7IJYNOIhN8wOBRvsuc4nrELWdV70
v0tTqCIiFq0BwPEzvxHEZxddWeDRyrHBkrn+phjHfSPJoyn4IpLPXpMvRKh55czq+rtrBl1s5eiz
CPetgvbJOpUzyVaDde1EfphteC6TtXCY1yCsmIESd8duf/4VqvBKPjuhV5nJHZxoiumjTUFq3fn6
17NJI9LPC9cOh2d2vJ266B1utnfRQr+3BJscW2+x6xzEKNmOrMxJB2qITW/80GbkoRqLzHRYICpD
PATYsUlyadK05XAWjXbPEgEgVTizOGaMSrO4HiU9FfCHEfvOaih0AR5CpPeetme2ruFejxt70zRu
ukOV7zaMxs/vqqFd9elc+mAFvdSZpofuPIdjfuecoUD0IKStZxsIVIaarh9nCE49YzJivumaq3/8
IZ969EqRROWPHsXRZqQrwVl/BiJo2Nx64ncxi5Tz4+xS/y+zwJKNIEkedjHv1UxBo4uauQ1p8XIm
PGRLPkBli7rW/2+hZEaoJXuYcHzxqKT5rJMAhzPXKipJnGxe1s+4dChFsIr8ZgDyMrWaaiyWi0cI
8dJxyzxcaXtkPh213G1irgDTDKrWgvBP9qz7qMj/Y4p8UdaT6BUJoAV2AUG+4Mum7tIO8ZGzQSab
e6SY4GH3A/F7Udqzs54GfFqvluidtQHlcrvzelOWNBmlUxSz61izeBVu1X/urwbjbrcBRAFnF1BD
8t8YDn5Gww70Y2bkf7pyPhMy9ILTCAVfibgbGBDhZ1NKlMVwXnWZ8f90ULyL7wwOg7oN6LVSSU/u
lfMidjKZe1N6X8i+OCddEsyPaCMeH8gWQXbKanVxeQsImB2ol3btjzbrbJZsO18uj7V469LTIpZU
SKOhw1XMjLcPv82Vc8MyZnkK/b1LGCbK4mkNaqylkllkdiQgZzYumXR1IsflpfVmZqoW+uGkXu5Q
cWNtPmZU24JFhwYeNdR2rtlz3mKIrQMNdmoYyhNfH9CSPOVmsD748s+VaFPd/j/4RsvRn8C8vSp9
tgVvDm8LlxNVg1jr0weQEu9IuOLLTQBWf3CCw3QxJiImbLl+OD0oWSxzvDf+z/nT3tmdnxGPgVxE
ca4tGw8n2JXJ3ptSVIV3+szKHIdLDBqorC0Uk5g36VALpvYFMFS/qkFFVpNKm0xgih7zbeajwcrP
b482Or+rdxZ2d2FHp3jleE/qfYHWLTwh6coYH/s/WjvhfNhzmeBFzoCxRA7PlLS11FEsM+gQbjK4
qwsbigto3Yjp64XnMhYyyB56qu6GCYgIneWfNHCak88b/nFgaHIpVhLhHDtvBdcWKd/4iynsPEUP
9Bmqc89E0dFJZsMcoXnA+B3dO8VTY4YmrHHijTCurtFLUsHjmm68jb/Fy1Rqk2ciJlfidJmkhtDW
4zV/Ewcq245T+nsnp7prb+4T0FUd3bKzWgrY53EEYUdo583ijPHXtA5D4t03LIW3QYN+gK2o0InT
4UmWzGm5uCkQrxbJVLWABeK4fGzJGw9/T5qSRii9x3IcMrdOpdKsSVo1jMkDDw9qjn1QGzJk4NQ+
DVg5TRg9HNGRxNqmTLD1JhGeFwo3tZmzVGlfnkYI0CDJkhuiKZ4VwaCKcJz4X6OA/obVkAZwsdA3
I1QBtRLtU+Cu6r/saaP2mSIjCZmW5eVTeBThC880OelxkNhWiowUZMdrgbN+eoul9tBrcyln4zy3
4hn1PXzRJLWrrkAMrfiwgXpQMgnJOLAkBDzSNs2qhUsovkdaAtcjcSF/KpqXlK0/BjhkAvufoV9i
Pok66U5fs1mU/ogZCCQZwhXz623O9Y46IxCF/DJNZKxRZKApp/gGqlB8S+nmhK1u3GyFAaBMSQMk
DoiDa1puyywjKCehgady79q/C+MeQbQN2y3boM8iOG0QKiFMMBConlnKKgP19+J5RStwd/7dCGIP
fKuq9TwVBlrhJUUawkiEcUDxQCLh3q5kNdk+LOFEE3C5tc0ApY+feKPUNOpHDDmzWhD8vXtBmADF
QuYW5LQBuzvvoxnrUxTeHVF2C0uAR01B4mNZixIGYBxbs31tulokXh7lKKlziv2VUsiy5L3u8Lyl
HIZnshHbQ1uU58ZVa2v+y/vKs9R+a1gliTz5vFmY4/FR7/4sF0zkq6i/n1V6wwlOVOtOWio/+/vF
mYw0k/yOqXbrdFLDmt3fWnfAv58mwv6+7z3p7+glYzj2qYXe36Z16l98YNsoAh6g1WWb2R268qxs
BvLHKwYGzD0pE3zIFCaXcikhGoGPe70I6aAkadWvImdrM15j9rXweAWAwGNxTdcG+FZMTRb3F/Nr
wyFgTJ9hdnsqHd6WEYHjWeWhSPZ/WajpOY798fRR0RDQginQyrtyY9+t2WjipFqdd7+xk8EpA15i
j6d0+G4yk+YHG/NsJyZMf7Pt1ileciUxjSohna3b2j0r3DIopvKUg14NjFVSZXeNbTjJ9cVqlQdA
aET3CH5dnUHhFApNRX4OpegwOme65U3By3BVE0rd80vtGhXAmz7Yna+VRtFOY0oRp3vX/EKy5v5/
SCHB5zY4dZnQp9TrzXpFpVarhyfPnfvP/opZIG/uNu2dFnaOV7gqjgVJKcgUQnwZR+lPFwsqKeLW
NbgLO5dnHFoZdJWL7C1wKsN5FPceDIlXps758bZ4fBm6CcO5koLf5IJjSEWK4udMnLjq+hi/65g3
puHLxgQcO53h6XRSf56cmGIZalHuk5PyKqRTLYbykCVAh97lsLLiXLT96QzngbX4swCKeaq7DdGU
X8f0wuyXjQkwhPduuth690d3Tgysvip3H+JPYuF7oT2rOFZ8zfIYYeoaAtxJvtYZRFX6kbtDwF0z
+4ESeN3RqYsNRAKpLpm9PUAsuWPDByBFULI66UmZ8qXkjy5wXAqjMSexB64I+LIjfLTUdeKazphV
M/j9mJS08FfYnRXU2kCaK0LPOPptFZRlfGPYk2a4oS9jB4OHZxNxTU8b3ZQNNuz6hhVy9YK3+j46
+0iXXPgKblZ46GpFyquHqXNjg/VMibwsSDZHgKdDpirfEummCpTOXgToTjuImDF+aqifCWs6SBm4
tF6AH3r3oyUTPYY03HwYtEzRTddkg56tfwWhUaMZuBUpP3EwyYm7FyU257tJeK0zFbB+Kqxc9dW/
krTaLETxAAQLG7DD3azCKtcbSE158wiSdk1KGuPQt3WqEcrI+bifyF0CU0nHpyibx4fC8qFcMGZH
EkXaO/hWAsfKr8tjGEXmiE9OfuhJ5cq2rHnFdPyeRJL8IgJYH61IC8NNI4pcP5pYOSK1lWtzgkky
jd9BcLcV/szvk9+FIJBj+uGQiEU1kcd5cPeaoTmsfkkhNQ4s95BxTH1bhwiJB4q7n98bRS+fzLJp
uk5BAqwVyIyS+StHRcVaWD2jcdYD32G/1vsW8mZYxcKc0dPHxXHhhX1bf4INWx67pIU/ixn8ktMu
bthkXFETCfwZp7/kg2gzc8+ZjIsyp0bdG9xMO9j4O7/wU/CULXcmsHkz7bW8VnG6LklZ3wOQVpwu
5JFSADXEhRB9VZRx6hTmJN12HM/kjiWYYsDkW05TUSODJn3sig7pSo+ofq1QFFcr3q304irZJim3
RVwTAw1UntZfmAF67X5zf4aLXbGMmMh6m1fmG582LnT3u5WnKQXTlXVNTJsvfvjd/X2UMbo7EYKp
ri/rQf5uqkKx3nP3e1FGVOSeb8frFIj/o8IUoGCeuI8we3lFOhth9JupVxsg5GTqZptkj4+RRNG2
97lw9cyPtgk9nO/r8DfP8x8sTzdJycquHuqz8P0rmoliJVO/u02T9vKiZyZWLJXmRJm5AvoO4YHh
8zt1LxfgXedtdnOeuumBEE90j3K6LDKkd7JiiE5ZKTbUSLdHEzMYRg7SV6vwKCUS9s98mpmy/MYO
JyIdxKD4P+AT68i3Bm3y2ygHHK8QWMLDoIIWKlEVU5NXAxbOkcFW1+HGjsqZrwIjfRsaiAmFvn9A
BOewwe3QOU4w0Wf4xAjzUTta/33b8DG2/qvN3vj2X1Gk+vjJ6h+ahL8H244kiLZ9LxA1dcy5pic9
qc1r5yAJjXLhlvUc1Z+l4llEziih6uXXRa/LR0yu1GWSzaqalvgHXXGnV0Ukz2jrGKNFIe3XiW2l
a+F/BwUBJGnhbwhPiVY/5Pq7KzpCZgsDSmL6ZpTmi3cd066WtHHJpohXYHxYyNUHd14OuxYofP3E
sFo5cDIsBVcr2Bn1qfsqFygLrP+JUTMm2U3UcGfL1AbqO32FY2TXO+oQkk1idkouqJfRQP+BsXOx
hWkjY8ZiRrQ0EmD39DKfKt2m6WJxtN/xAwCJackvAAPzwwWWGXqzGUnU8+NrrXpH0qgWwyhf8bDe
77LP/YdYVUE8Q59LsD82pDlXlc2QnNuy1YAEI9YCi7XYwylB8stHP4END5NzAlkxOSMTW0yWYGAP
syhHxVvm3YDTyYEGmOJs4R9cfG5+uWOurGKbuQ+RRaZhNyLoYIue7J7jLukwQaKw2QhZdJWFGFuF
NiuRqynSHov2Clg6X1R0U7J49rPc3CVfSpjgO1CyXN6pE9ZTccTXgFtDLMFCY/6dR3uqFm2UdTqP
gX8myqmejuLP0szTwWbG5liJkpo5vz4NLll2/4iSFsqcCcqH6mkGTpqSx4gqylB3H47MB6RgIQiy
Y6LtzYopX/sO4E+J54Mk49shpZGhjhW2b8xM+rrm0iQildL/WYnMD+gc22m4gFtAic72XuFQet8L
hLDHV94VLo6CtBTF6b4UJi8zhNCWBBj/0Kpg15zCvpysHc7azWiSSV2B1n7uz8VbhlrvUkT51hC9
PU6NYf0MmpBBhCeOOJeG2jouZYpa6gMxGmR0Byfgi11Jen6lrjep+PRcxxURXiujB4ditHaZQEsK
tAQnPlrTwsAAl8fX5pthnEZ1ZVpZE+wyGJEL/fSEp9jiG+RVEIEI3LL0gAcqGYzG3Hkw8F3up8wX
EocphEdhR/ROZxmiOr6T4XcpXKuNdNgKgTi4wd+he78UXuLjx1Kq5BOMStOPODpxhoPLDVnn6Qpt
KJmh9k3B2YG5KHtbcrxO5VCXqHc1rDN459GqTEQBo/VhO/W7LL2x0c1WHMawec30DfIEDjdYNCJu
q3yM3uSB0cofaef6oFXfMSuPrALi0gRRMGdlwcVqwvcUJOv0fUC/3nblwjtlkYH/3s40bJ+QATUu
hWmA8I8I/DNbaFb5435YoERiqu3O/byZdMp1Mio5UVbiLPN2807h62n8okXG0nWpbn1tBUhmMN+H
5qj5cSukQMkpMdiabmWutaKhySz/AfcgvTbrXrULgnErGHmnillEXFhRPO6xIpEq2As+ypejvSVH
6wNDUS18ANd6Yhh3CP7Ig1XUY6YOG/JN2IaVQOMjt36ClmmGSkzCmKMP8jOmwQsFHOV8jgVIPaBK
ZOf0mE+vmEKtWv+nT91fvhbvsCJ2xBxVNeYTbk7L9foMk56vUcz0lIKTBSHFMyjBHEf6naFhZCc+
L04G0FQBiS5Ukmzg1U2DDgzvSvLFFPBevT6eZ+xVFh2lv6ldyYUx8dyeggjFsOeicg3weOKjP0zc
6vtXQI2VV1t15GQwu1Xg/EBA2bPLW1JvWhGD8uiPFzNtV76kGDk/Jr9ysIJan7JhrmXJvBc995af
YfoYr2MRog2VSCxAZXQfw4r36nQ3DIHCrAUS5GTFfB1qwhToNzQVEEXKcNR1MP2dQzy5V6IAvPgo
2ElFpd5DweA8Bb76/w6Pm6TYvBD2Sltup3JyCxuMw1KfmMoH4lKkc9/Nir3pwq3l/i2w6xm9Q27c
LA8yHEUVuOSJ5vbr0zEC8B1U3nbAFi7m53g2TWf/SetMbJWbdjpMcfGMh8Av2JeU9grica0U/d7g
LLBpuZE6WWyNTR+8kiTUTtoGg80FTvEsJ6FNrQkzRN7QJwk2Kw4PzOUg9CV6QJnioF9RIsVAWGZx
fj107yFp7mwS5nZBMmLoHT624ZThCOGS+NsHHonJbszF3ROp5pqCOHAW6dapxbaZAHhTn8Qlp00M
lQRk8dbSqmEAaYgDKHljHjf6jiFkGNl9sJJOGmKFh/PwUIeNfW0A4fDkhYeDZip+xlqCrwDCqOdJ
7PLaGtgXCiiXyRAUv3bDbIXRpV3b/cJ9vD5XS7n3rZhnIQT7PDWmHn3nqL2nEjXi0lqfAH56bhXj
F+bLnjhfGkGEsCeOF0WuKDrLhEo5YJOLgSrWnu0tt1mr1C/WzYe7Ssx2KnXpIgOOqd5yZXbbTy62
SWdtwaeoHxAN1N0F1CPu9Ikg3FcmPYq1y7PDqiyeZArIn0fHuGlpOh3OpYj938dgUUSSaICEfcKS
Xayqt52LJpChbNinVuxHBOzdTYL8IGMEA4FmLYDwRVczKhfeg/QDOXI8dKAHhg7YrtE0ggHcMw9E
S+JTafFAWNHPvhDgJOIoTj8HbS8VMDnhhYUwQx+XTRg0gjX2QQ11/c75vD5nVvI0WhN1eiw1/nYw
B6La/41oN0YGnkLwvk5rSyBnordgPfxTgIg4WTXlW02Sl496Ivz07hujjjmt0s1muv+OKrbkch5x
tE7KWu2ZS3Z3FSukfIG8+9zIae6ejFvDIoRafWRFkpjyf13nH6A+v/Bb3j/MxFATVk8HtfXWnWBz
i47R+9nh0gFss7XCMOj+Du3MFixaHeehO+Rs5048B/iTLb2kJ2F8EmQhWlWGiE8WF/NGdqhwh56C
TzIviHo9oYmwt5mltiep2HTAF0LvRV+JgmDIumrJmhCw21L7G4o2Jv1WlrEG9svUh0h/YGaSOxBq
WbOfhYjVL7YmzZhaAiBH7ZLAVvI/zQvl4X0KGvp9m8eIo1wA/9chfNmO3nad/k3AiAoc3q0yLhbk
xVlgd46vboFyBJ6ChwhLg5rRXH3GMq/c+5BveJ94jrrcPRX1o4ZEx8BIOzsA8qnI4GcXPeS2RWqf
xR0z/NYqPTQDknY1O2aP/cHR/sCU9UJ6uvuyKNoe9yacPM4XFqhyYn5n/svEbZQJgCKuQi/gtPxd
va9ldgW5pW1+UotQWhy2281k44GvZ4RrKEzmtEXUpTHO9BiQv1S9kckWK+pvMU6tmkbm5/spMpT1
r1R/ACjiFBvWXxAgGqDfXpax0tEY1HB5mjgIjwt24BjQarzwNc/fEjKsUiCIW4paO4UTlmiMP2/Z
Hp8nS1GnuUuB5CUDAQKUZAB+Yp3Fowm+lThquPIhxwGB0kV8neLc8fyuOObszMncK/39FAVn2f6G
BMSujFpmuJtpIxMykBv6IBLlFU3dU2HZ9nTWYnEl1s4Mvb3k/IsPh04ksmpSXh5BK4Haxjw4bHVE
yx6ne01S2OduKMm53s4oCyh4Tw3WjcH4o40gg6zRkVRTyxRPqY1dCZwI8+Uckla0616vul3JDqEp
CPtmsZTbmewF7TNcJC90l3QXuQsnCeqxV2frOTJcgrxDLwxQpyyglSlzejd8TXqGyn8yEf1CXEy3
fBdrhHWgprJahfOtXefuMz23ZThV71i2u89ssbwh0tfi0pYJ41XyLO799KzHtKnHSZie00HJKur+
u+ku4vUueHuSiI6mozlSGBHD+JYK24DyEepgtHB/q3Sb1V+pYSGe29VRI/T48JVrOI8jJSnk335V
CFld29uHu4vPKMwbxChLRqQBGTi7vGYP5/jgD3uuw2Ju/Ov4XCxK3LIuMBkXFgz6+tZpHhDxIPwm
kSlrVhu8P3RLI9ltQVxBc+CR2Ld/fllLdtEznIE+My01PpgPfltiw4dP84dnE7BgClUdrCYwOArG
JvCdCcrN/iRySPfN5ZEQMm6bfryfWNMQVhAslwtCHzhwR5Sk3hhOSP50i/2FaNBcHovbM/hcVqBF
P4rzWght9V0NG8qxPtri58r7Ehap6kOcIY0g1vEDVli5s3pU4bjMdot8x76yMqcpUSHsJi6u+CxI
MeHJ90pJqUmz/vf0cWR5vcNpSgh9ppj/ykWDRYmCAjF8qAXTyyeio85ag9V+qGoFBsthhLbgpiHU
Q5R7i9TBr0+RoKAl1FWjLbaOYdYLz/BJs2p//hjyBS/Woh4kcmiLHr6Q9x9/WMUv2i0klyXsXngF
e9+xkWcrV8jsmriq4Mn/F0YYQ7U7s4vhRcWFZQsQLChUd1FFFAxK94h516W4zGBbCGhtH7rxagFh
rGSYzhEApmmtKW/eWIH+wGCVkZP4hG5BvJ8PuOtLCkxeT3iUNjMbMpvss1LTJ5y7nQrMIKq0Dhjo
35nUYrX6/cHZ9eAMffpHxhj47lSEko6ZIC/9y0TbKihViU/o5CHc2BiAaxtldyzed+Dpe2Hg/ptx
kqsLA4F7Vu/5JKnbtqRdZIYO5cHY8tm65to0omUkCzD84ncBGPsBLfmrZDl+vyFNluM0Vg0F3IrN
hFI8BtLiN2Q+1LRNdyyPhKRU0gLTLyR3YLe95+PIC6zZBvicmwAvQnTMAGsckhdt082Tec6/Nlvl
THs2CBGVBQMCOLfHnN4qlei45KJM1IT6p43wbAsOnwonfrz12+BpBR6F9CJtUdRf3sksEbfyFesC
WpjS/ITRy046Ua3gC8kZ1UcTtPBKW1O/BH3VDI0+kjir1/9ad7PPHZuKs0xx6UKiaBjGa4ghZbu9
tvPMQHZmL+PS3QgJnHVwZqipDuEfty2bIBC+oZgeVrGyWqoKDTBSpzTvc/uTEyYZUsQAdVj7v9Lv
SvuK6i697GjazPIn3qfUPixep2erEqr6S41FtoxNaWtW0QOPL8x1cVqNZpT2WLrSPhaFnhgs4+TP
3wzOTohwziYGOKC5gRzCdABeIM1vfGZN7jTPS8c5P0ogMw1/iLtK3kP57mam2GABqYs/Hna93GGM
5Wa/A+bBKrxoSzqJjsizORpK6zWp3NOfFvSoed4gLNffNFaUYniaA5RRQDYbKnK2TnFocQrk0vtB
Us0T1Fn72huVS/lIJNiALCi+s2xORX+iefwBqzUXOM+y1pxCAYXXs5Tnsln1NreEUvlt/L0eqeGi
elr2cLX/wJQRXpQBSxaBstyRvGXRoObYAo6yyzR+b9gmIZyjD899qGmM/f4rlKg4emmn+9KtdMKx
29k2r8Hu2FJ5kHVQIabPGwYjMwD7eH8t+lbbTu7f7adZ8Gj0pUNai0HNw1+FbrvQtBJS3BKn6Jpr
/DLtbge1zXD74vYF1kqrDTjSBWlayxI0Jl3F2d0y6N+VA7dESH2syb3OzJHOgYQ1OM5vqsE8uHB7
y9k3WSpEo+vXmKXbiSW4nMVN4EdmZRJkWtT6+jmgnPXJOldG7t571S2cR1XxA9+YWf2k95S/7FCX
wQ0rmZBzujGly6xgKNvuX8HiVdZNVu93wI2E+D9x4qgkA4BLVLkmTHLSTKpXTgvmrCQO90sYrYk5
KxaCfsRKyoKyW5IIB4mkVdjGwxoLrgdgnNPZiHgYWhdwTQsfnEU/cNHw8GWrxskBH85f5F1ljKMv
/q5DPUeHgUNETSGYVjJ5GgZ3tF7l/8nm6AM5cKYwh1a2yiFEvjlhHKhcHJ+nCh5TYVBwUFVrQbwp
BJM223/jXo9jznuwkPU+A+N8TPU2Ac/KYYYz9ApiFNEP9Ogg1npsSmoIQKfoHFbaKJo8N73MJVO+
FcKKiejYz+H1/DjzWdX3IDhpvA7Llh+bfWf3bEWBqrW5xxGvSPWYPdsQ7LijrUqfXKvPrp8M3xlT
SMVsKlCNDybHI8Ktd9kTu51z+XHgtgw65gu5DkbeHtXdZG55hOzf0Blq0m40Cl6db/1uEbz66iR1
E1C20VlLrtvwt9KWWSeXCjX+lQ5MkyjvnQr5T6/LhxyurNChrT1k0R0PQ33bnmGDLzQVGokNC7Sa
ca82yx9k1Ly3ICychKWX8WABPagoWZfuE0MFAI7v3GbeYIRwJsu5yg7ghTWIFc2rlhqal3zJdww0
SDUrGzIQXY30Ynpmv7mpoIXOdSvT3d8vjI01IqKDF0hPQq9iJdHZQbx5PcOwooaqwITdUHvgnnOq
GYS0ZPVYx7Gh53rBsulskr4N2TgcKB0wJS4ih99PwY8HY1T5WXHX1tXffiWy29cGNfjq5HQi9033
ZSFIu18xwz3A1ESOfBq79CTZoHbh/SliFDhECOMExis5brmO8X8HYVBJrofkNvSvISfUzP6zW+yX
0urR+gFZD4kXYDXEertj7OyBTbyZCjiWspn7lnRkE8YQ+UjVmZcLjjesdlx/CZHDnqq51UD9I/Nu
otDxpgznjH6beklPPMPePm3LY4UYdW1dchQQrVF4cEHQCT4upp+IfGDQMK3k0o6JkKzJOdragxv1
rrK0OdtRDNTwl913QWc7BOkkx7R6LIRdeVhZDmvmy28DK6zvmmg8HQzmENkfgvRCRJziV55Ni6M/
XUTradB/6ijWjtSQmYWJMg+hjmSUBd/6eULTin1QauEM5wCamIU1uKt/AzK0CNgEzoFBATAivAVr
vEWJe+dGjPXfNRrsOjhfw58R59A4mZqy4f8XXXZyg/zdYQm29PwEzG5TSfJpTEbaeYiHZxjgFo8t
QsOCOO38KBOm6QrJeJhof3W8sms5B38dbrsdyY1VyOyboHDt34ti6HWeeTEe/f66wyM7W+GM42Sq
InWLl6VnEjKLSYDMLp/3eeYrAOjv+TVEVUDSJFE2gRksLonNyZY125vIvkRA0eEpVMH0bV2VHgMJ
z48C7aqH+xduIHgh5B11krlCW+Yry5vSZUIRu1t1+mZIuzb7eCTSyRfOijk7HcgzuYEp/s3EKvUx
pzjZlDpOpug8wYwzKKkiQG/0omGBeHlKK0PsOyNqpPor6+hEHMJbhBWWFlboQAXiaZirsbFj7pgx
ZT+QhSFcj1JaF9PJG+xxC4nwjnE5jY6AMo0Y8NAnyfMic2iVa56IT6OF5rjdwHNuLBom/ozXMt2E
WZOw3FeruKOR1VFMg+M2S2rNeSf76qsCwp9j+hk4/Fzmknev+xUUj7tUDtBqFo217RbFzm0igCfp
cf8Ugxw5BUa7dWUpdnzWsE6Y6mkPb77+3yNUQ7+v9HCQWmzQY6nj+BuDyWsp7nx26RQXwU4wvADk
gla8cKIeIsgdRmXGxQq4F4R0b2u8MHZnu25Ra6RAxtss2oia4W6sL1IW3egSZ16tAAB6llarYpsP
VBvWUy+C8W2erD1nMOk+2c2XB1VgpWi4bRqebw4PTBaFPZanquTtxuqgrEBhP7FyeutoJsY8WG+N
Jzuq8Js612TXd3VTNf9MQEfR9yzq9OepTKy0HaIOix4A/yzKKbhLtbN4PhqlDQe44jBLND1EYfOl
au73+MdbG2QA048IVyuyruZwjfBFMSZ58tdafKMYAdOvOHlUMdj8BsSbwAJF8wxHFaXtqIr/yUrG
cL5u8WaYO/Y5WomAH1I0hRPu4gyxyUaiVS8kHdQeVUeldHLr1imXvv5T5YKdO174wJ7GaSqqQkX0
0lG7Awtf1AT8zA64RY4sC4B/iS0Emxyc8fV6SR8QaQ6HfnO3RJVdDPtpUxxdcrXTOf6Iah2x8blG
pMef8Fs8rsZxBEXJvE6wxPC5O3HXPuq4kxcZLNGAsSVAwzcBZzNo8yQNV06kObfDE2tg8qZ9kRyF
+J91ukRJDCmEI3JeuBgzARw+32Obi/Saiha+y2IjzQXOc70y5upeM5ASQq8lGHBsQ7QcQAQ8tIK+
SQJugrtlSRJYhYsMAi41X9axonB7lAHWUeCNAFGWuIWcez6AAnaSJefln3eQOaYbK1klSmWBlwvk
UjVND1tHQMl9o00CMTcq7RZl/npOPQ4XtU60Hyr8g5LSSPIXTs/2jwPnf5JY2jFSc9RUEe4YFH6v
iZESGRG1trCwyZ0XcpYs6HMuuk2W4BA3cSIR63GNNEtPbdqxIqdZn4K/7PZeV8Jca9L05AQGxjub
V9W0GZDeewH7hopVCoJDo3DZYlswFhYPLwwNetl9llRmfCtpD6lmP/Eu/2xLJO7ToXuqKXoPCF24
euoFBKBfJdVfjpsxIR+uJ2EAZiyHN6rNFKu7ghmJikt/w6dLNqcxWafOnZukPB0CUZjcZtCCmERy
BWyxFDp1KLplKEgRX416DKa3v5o/NnNlh6FXN4vFqf4bf3gc1UxIxVtVU89xfpxUYXdzXYClQoEK
5lJ209UAXQtxWNN6Elfee17be7bCbKbPtEE0Y+vizd16CrsNqFspo3I2jGIoizaUs6TZNFQFqfuO
++zK9M/5Hu+GK4zj7VX+QhkhFQErbAslDwGrjtkoEbOyo1/h+98VxZBt88tDvv+i8KdHuuUiH0Aq
DeaRJ/cA5pJKP/8Bz0X1UEjd9w6pI5RBzW+nzyUbK3rTujK3WbrXmKPP2h/b9y94OQvdP72Sq2Mr
UXqUE+zmV5HB7t6TFK+YUQynQxbRlfEEbJZ56Xp+JzCMwbcUD7pkYiOW7c7HEUEJtjEK2ZNSunHg
XN3+6lYtw7uM8ylUXtc4yvKJfYKkKxbKQvcvjIdftzJVTuBgo1MYJPMCg0Gtl72xHOj9gY/M455u
8YocsJcAf0r0T3cHj/oilQuBuiT91bxZ1ui3nUDL9aKTu/fW++RbB5M70M7sEHFf32FLBjSzv+cX
lGio8ipwUI4nr1znuOBbQaQEclkbJopOzJ9Aj2SVzhZqAXsc8g5G/zmAz/y5+0Zl/n0rM9Tsd2G7
PRBNTiYAUzHgJolvDzhvsg28km+33og1F23vjQcw7jqDarOP2xwVALhhMbpl6l/NtdilIomsFc6u
Zcm7CcufiRSPwQxHrPmswNjLR93qEhmgFxO617GLTyGPQ/HTkIHTsqgnAieOwHMsNSh8t5IXOGa7
smhh7oQLo5o0N/aFxepBdZu/RnP48cNTReY1cA3ZHuuElC+bChwdFtBnGd8LAqKs0CAsojPS86GJ
NZc8VKplvLuhGgkjzXA+vB9NI2jNMSYjirIPyA5lRqFzrhCZ+yAAEIuHKVk2UZaZLXj9qoWRQERH
5IzradFh7MFHNXsbEGbQjNaqY84BKltaQMbBrd/24U3s0a7hfs91CZLz/CQbaa+dlp8IO0ivk3q9
lgq683kbB6bPPcgV96WHLU8qeZkXxrFOWL3G8WtOpzDzk9JzRO9M7UgJXHyda2ug80QVe/J6SNeU
UVbIZIiPegHpSeL95kTwG3qTL9nl9QH4g8zOp5AtioGVxzdJrhuBfNlDrN3mzgwTrHrcnmmMJA4A
DNHdky3YewroADUaFAcZjBO1GaRsmvjkodgEu4fuPguEKK8avwHiv3Rohqm330UMVlh1zOUgX5gq
uYVHJJyauwrbvypBj+byc0T28efL/RQB1MbvWCwNyPRGpYMH8zEOOYL6TaC3ZIiE7Tn9SSiwZJkg
hJmtcJIH5FfNf8r+x4vWf60CoC+oZfTEGG9+odNr3oxXPyvj55dK/FiDNWULoZ3YmN/ku1T7APc2
ACYd51UydBInXQYrkdPfC2uekUvEuxqJ9VFONb9uzeJXF5BwIJkqD35cSvE0MJJ7O6r6UGpgTtyO
2PbZqt6YryazkbcF/GTxb/FBC81JRWI1PeQBOxEIdUbhf1P8icHDL3SpKFr/j5YSc2ZCIDL5RM8m
RRJx0NHwHirC3bG7M2HkiLbFhHLDTpUW4RyfjSXnJTgWySSS0eUG2gQjegxeTI2mvRvV43damEvJ
82708DzGLGWf/XIYj7nz58SB5I+Y9TtJ9ijfvlD1d9gAb+iIhSb16Bhrbb8rx2UXN1XD85/xQahR
Mtx7qikuJVX9rlnAbcxmGBUD+BB1u65DD7DOyrJjwshQg5vPmpYvjV8xtcLJRAL1Zm+2BhrLEHfc
8ixTzdcXoyvrvLTJjUsspf0kWpKO0jQ7TaAGaCLyXnHHFXR/dWZvW/9SwFwsoy+XqVmh9o4oH76k
FdiQBLwvG7FwZc25ae5kxn/rnMWh4Weas94zxJu6KKINscE1iHX9dCK651Gm1+3wQipPAccNLQz2
chT3eOpBNU55KFC7SxzFt+uZgqb/P3FNYtlxV1QspFPnPhQWfdGGh8jzltkEdYRHo0CppsrRxhqv
GAkiZY0qUeRMU36kQiUhhZRV8gBVF5ZWqvBoTDm7R+PvN9+GY26OaG8ITUcN3fJYJLJTkZ+ZVP4+
zn6MP6/I+FalDrIpX1jyvmFA7NEm3pyvzKu3p/xbrmpSnPU43CH3fL4BQ6N5rHM2fmEnwqf6t+8t
u1XsGgWxEEAPp1ShZUMCGhBkAlK1W2GEOYqRZqxPDD4wDIb4DDOoK3NZeJdnK1gMEf7mhICYphDm
vuI1TqO5l0t41JBsEulzTviIMBwMW6adt3DH1zCzshkLajcbQ6TtsWoe99Hk4mqM0tK3UQoCGWe+
eVukfNmf06oTGyZJopMHbr0MFhvLCSHBJUZn3RBIrXS5bpxW3m+JTmnEmhIkxvtBlnvmXiAwrmt1
R67xCfw8DqSh61piasJvkTQYx7gqDRlMm5yxhSMl20TLR5Ji5h2xiQUvfPAbVB0PaphUXOW11frG
IKi2M5TcXycImN+iEcL1quahwB9cv6KB4pCztupgnIr5rs/q6x5KXxwljBzMI0pXt4301E9qYOb2
ky1UygVReOpzwVPTEjyoF7qtzCitJG4t5IUAyUnQDnKtl5cTFdmYMOu1XKMseNMsohkNJozZ5j4a
uLCj9grXgxVc/JpbKmU9vvPVA7uV8iKngV5Yo1fPxMcHBJyAE5g0Tw3pN07X91+SlbAlI3LtVpFv
rexPo2ATODcs7/mEkjz6Yx1c/Ojav1tpzwXIb5E3HlHPFVoabgHFT6zeJmoRjFiFS1XrIFuh8fau
8TJn6AfipjT5/0Dnb4wkATe11O3puBaAP7LAF2wDPoJiYmbNEou8OQJ0BHO165ER3rEvttYaEn6c
jTcdPrRvzi8csXdOC/f+VZXOn5IBFqG+JxE/N91MyLy0aEQu+jbwM0FbzOIA48ZkdSHMVytJDXEo
X3ajhG734Zc4UpusPKW2HJSE0fHGTRzMUnaFecNLEtPggoOyFWQ6/eS+3BjkInHYis+TflGNOkeh
UCqCVebr12HEWM7NyIpZDL/MDtM63EvpDMhR14ursb9CYxDT9hhR4rxlj39Wa/91EyIqRNIPGrj4
lE6EbuB+nW5P0my6muA1G0auZ0E2WAnpAdFq0On6GrYUt4AquAmiPSJhQgGxF57wIekWnxxxV901
09w9ycHogsdVHpUjZwVOUudXLwpaseJN6QZDwuXXyAgrONMbFWhjF7yO1ajKss+QqGzKqhzuypIX
0a3yrwydCi/H3UuJIgCrCzq/7TgweP7WiS9J2HAa5ekKwVRKQuUfxGzIOVxHikwUFPuhQqq49jwQ
d1C0UmyCFNKit5Wq2Ag4ykMyNOhorb2zUtadOzcy7idiXkL8SCzXL4L2uc+Pb5HeAcC8e8Iq3Vnt
JRPV3/oUUlwvJHyZDy0sMP2IiM6fOgF+MHCYdio0f87vwq1UsLs6da/3gRVy+PbwF9nfoz95JVTH
BNcfc8THqwHCGRCt67EnZ8KLaw1lr4phGBfCyI+JnMqmpXpc/6QmUAwDnXJZPWgB/0N+B7ZRG6oP
iwUMjv7kP3ZknynnZqYNZr3ZmMFle4iG+IoKNDWUiljAfThevM2YY+CU6XzTKXrhxqBc+4dYQ3IP
eIdAnBl8weK6jIDZDiT59vq1oBJY29TXRDy5SPLDkn7v44Eqypw4KAUxGTBFKLjSKFjZWGQacqXA
w72ZQHYt4N1eEmrdsd5xFONcQ0XogVoye3HNccDxRNrPMDo4IJdb6Y/X0ay7YIhBOBgr0R5UA0zp
wr/Vz6HQ0yd6e8ZzjmLCJ3TsWxQWq0vJ65gABTrqzv7O1T/Ox//kkGqH+FcxY6qJPFYLGVZup9VE
jlp7RbDtDp7VUkvwMeI4hdESOGPn/3/v92eNA0gFUsqpVthWIjw/SAG5RCtdTFzhPMzA/kYP7x6a
3T8PDDoLWn7d2rlcGbFlpplzckLQ5CwZFSU28cAigR2lYurxjwi6mm3tWTxXB4oDRNHuJN1ZLjZ0
D00zmhKupmrQVDu+T5MgKeTTmKDYiQJdeYQ/VPJYU0h6RYOoNNIibaEqesGd1+ITiPZYG/w9zllF
viXsVXzuShZP2W2TXK4bexbToufTIZcy1rJNGoExitt7z/REDtZqDzJp0jjPfS7ksr+OTby4xH8z
ozM50XNLwgZRxDeJPED/DxGYqGW67c6km1flnWCt/QeU5zDOv9EjnAvmXbuamnjfu/4m0Cy/Zuq+
bzUl8iT4/SSXoOJ7bFYN1ehYstfUThcBCoulHO5ubcJyt/jcYkHMutFpQlMqosUEaNCnDFlw7426
s+ccwzlN3x8a/hxjcBcpQLI8Q4qL+JwkXh0b/YRN3Pgc7A5YqP4rkDE2WtrL55AoXnISCF2Zvd4a
XUTliflOYiHD7kpXYQvijfPg9Jdh7KvzN+8cBXgeju/W6NtvdDkMDsbfMivwzUVZJzvpgbE3xG9f
KxIBpNXb/jhafJEZZsTXI860wreols3f3pctXAndpustdSTt8VS5st5prGPzaZIo4JlwBhgZ39Kp
nHBYRlwNFqnvOUkRE6bXxmydxj/82bzCluyVqQzGBGwmmtX2fEpwPtLrfvjc4YIROZNmmSxAVJcw
qnOBIza5VQy0GSxMG3j5TkNOcTfknAGVIo7o0k87/yfXN1cd68OqnsivzRnMYt8Ne+EsBwKE5TwC
BYxMRUy4KR6g82n3DkxR3q2jMR5ka3Hyzg2YKRQeWxABfKk4+FTTD58IJY34mYHII1QeMyGY8mF7
VdGmhdeG92qR+tAMOtRCnsPId1VFdiv/jUDdKcbcdxBQsvDuWlwYwW6YNGSMAJxbBpYvzfcSfHgc
higZb+KXBPjEYoO9v4gCO3jHGH/kzl+TZnisL13uIlkegxGNf/iTGhiKY8UBgezGaLAsnxuTqr8a
nK0xXP2NFe3hg6yyUbd9Bty7maBYFJP4mRI3UfpPuvHI+zVIurjpu66S/MloxWKVgbMWOZK91aau
aRxLJ5XAQy2w2v2TN7jxcDGCL01YVQVr3satTiFE0jPMPJb2dEJ4oQEpXa53HrgTLrAQJar3e9qK
nzyBYZ86KmjggRvy8jtbfLV4Y760mOW/VubQhjvBBACri9u3akGxm03V1DE3SzCjTEIDcQsqe2xV
a+tG5mZmbo+3JYPP8qzF4x5IoGh8zAckyMhueJRQWF2DTI5gFZuozFktKL7ZJ/La2978CW+f5tcb
pHackGVeevMaFSYcPqS09bZq3SJhTs+J1ZDBlB7ig5dUkgHQ/AOyq0vzBVgTmM+ow4uxxnK4RJkD
3OJ0KXDeUxRH0CTa3I7t2n5NmMNt34bL/TkrCIaCIancsVsl2sxM/pVrQL83ofwYL01ap0WazzXz
xkzuBopCOkgal0TRq0Glx0evL9NmeSLx33A/y7qGrBst23mkw/z4yWtf4z0ZuvZBhpZx1wWsbGqO
OqwXqspgeJEvwr+20pWZUBidTIWiGnxLPwse6Xqb8b+mEJCCY7/lPN64PXG4z9moq8Xj/8Ub5Qoc
vx1Pxdwr6sv1TVZ5yX9hAa+BFgNRrSY+cO7Ow27Ckr0yQGmJa9P+1PvcjVWZB3BBEutEiNyN2o0c
UETg/MfwDisos+CliNVBpLagzNoOKA2gXfKR+n7aIk/D9UinV85NqQj6bC/PyfEvaKVjWZOag4zr
SYqjaMdwUGYkwnoQebWqAXul2FQZL1SwGLnJwQk3vzpJW557LEPSbFd2uhtOuSJ2AhrmJq6/N4qI
YsLY86FUw/LYLrMxDhpvikh6EHm2MeKM4pe0VNxF48WLx3eJc8smQTKZdUJ4KOFVsI8uqZGKhMAh
o7CpqTdijdZ0kZl8R4sNgU2O4Dyu2xTplSSzcT0s3MxDDpPjWB0Ie1UNPAuMXhcqphZ3eZSeBVVy
HYDWXDkLPRsgg0EQXr1+In8IRrSqPKfkdgn/cJm/lNYMAlJsiJBy3b0EQGLc50H28Zsxs0EaZt2U
/vuiYgFQ8SCZBV+CWmdgO48T1sTv/ZG3UviVxrw/UhT/zh8uPgnRucwPEpNJ5W1CvNED7/SHChBd
InbvGVPAGnOWSjpZVzwHFgzNDfrfj7GqFZufLJeAL2h4mgXvsQYE/1R2DkYvqGWKx7ZpYqMDiBYt
OwdPI/yw8VEHkvFa7VpXg3aQa34KaHi2J1fHERch50ucCNqerwLoqOT78AchOXPzS32eKkWW2/5J
qvelYr5KKAKopj16WogbPUsvvHGWAUgB0H42qvS6G2+UrP6s8oJn8mt4X7hkfJIqisLT1DhflP6Q
TQ364KbxNqa2xknNH949m0XsNdOj70B0awuVd2c4P0JVZOM1sV4B5GixH/l731RnY55bnp25qzzN
e9CDfZhZLBp3APB46QPN2oFD45oqukxHnpi/rh9DW63DHZQVnR9Y9DOswH7BqVaAUaEdUwpmnyAF
1nAAjMg1O8nfbHq1NUt9bQCXM20mJBnsxBj2g8jbySpPkWBij3Tq+DST2Nw1dbahyMy07AwHcI5j
dM0MREJOHx3UviEo/ubBEf/mPCX2439z5vSsmOFT/0rP+p8GNtGRHKdmRPYYAeDtb9/l3anUj5VR
cF1lc7IyMr0VjbDrkjhLXWAyMf+3q/SDi8q8p80VK9jtvb14wzXkjA+PYrl2+1Sg0QhJJRDM/hyd
59iCZESYVpz4oXqpSwrgkEQUSpJNsVRjUZzBdTwno8rUbzWrscLGCaqfpPIfiUVGLZS8aU874Ucp
mKiDd30MlRweq1fbd/iQR5AgPcdRhx29FRaoMik2+g6eKyj/T9rJtoL0a5YrwC0yPCpP4LpLA3vK
8nd/eLRBINGDKOmDVilFQUDPjTWWq11zOYKJ+faRA6omXbS7n9t9l916o8ckhkFhihekrFXd5Po2
mxyIAXDgoHLjiBrxsG2AMUTgbgv2NkZKoXW5DkmaOzMevj8HZrUiBRkYQ0Dw0kkYuvzsCVkWcYcG
MUd2qTcw5DbdIxZnY5t5neS7cGnpR7xHfJqLHhf2PZorejXu8Dzir5lI9zxOtBqnby3JTfk5/7QD
CKl9F+F5WlMtAhQm69SqHqLpoh092wm/Fk3O68lC3ee5lRhpCpWgKJbtSUK1exejPObifuD4g2v7
w/zo5R5gq4/aEWh7TLmdulA9cMpMa+17yDrpHGkZidiHKiCyxQ943JEPr0UPaJTONTgaDa+/6T18
dwSwtfOZRrkpwUMNcgslEeuMQFR1oF9VXmfiKf58H3GD3xushA9lGQ35hneu/TFL+YHes/3hSWaF
9WdZnS5tewSwxqGdQ1uUKQAowv+qGbNNi1Kk68CYRJVpQdDAlAn/ax5uS+G3gt3skbwdVLUuyLYF
u8XMxkHzaHw5IpMZijrkiBWi7/Ygtz1AUA9wpeno9EaAyLmjazKsHN6Sw0Nvrg9K5UnbukZvfs72
X7OnFsn1EO8oTxhcnLLQVvZW5Qj30YI/fcTExan2J41EhlUSRKj+FnYfePqGb8vjl9yTapcobvow
GaFP/B8h7l8wIPyO/3xNhV+6WRM5BlvsixiEkeAeEEx/LKwpBwOIH4pPhhA6+FWMHcgqk556sWPe
7Oc9eKjcj/7bdVDvOugKcYhGRksMOQbyAl5fK+QWFaC42S0cM6qAgmfUZVjh1nPDCFJcZVhcI3Y2
8CkBziJm2sds+UvbzkzwiuEdqtmSqUE394ryaLKAIx3Dt1kxwY3w/GPHhXYiTfrVDHdh9zbEWxLC
tk1BSKgMiMc5Iy5qgs95BqbAvC5nthxIIRA38TcWaPAMhX/rbbJxRp/9/DoG4Y1azQoMgilVyNm3
WZlDEehHA21Hdoym9D6MoislFMGOqPVCVScoM4gqPeK55w0QGh0deISaX1V0KLR+hr4W/E/M2hOR
pQBHfV9/Ap9Gbcjt9q7YfiMm557HFblk1SWDtESfNLVjXBwkOpMmnzmHxSu16GH82XAqkaXGrJeU
fWY1HmdP9Ax1XQj3yDGn+8vjx3AYMVy/0kT5OSXQL4T7meQdmhyRK/7jIlV0z3zFlgw1FkEuyaki
1Ig0OtUCNFSMY17QoT0twoUG0xKG8yKuvSxAPGkybkviSOe5BERVlaV8ZFqdt+EtWrq/+m6fOlJ+
lLrQRBu7YYot0GdWrVkGBawU8fOgw3Q3z5qKh5yX6UZ0kqJLQHGsySWjvh4lE7Z4yVloZtHJb8i3
P9aMIxkQUR8Mtt6qHcVzK3R7MTCRUzmeewqyi517Gqhl1gkOzWdJQYBUTpfaydN19cDy8ezd37w0
wgYiG+JsdWzVTmZH3M0rJ3fCG4j3ivnN57rArETtOe9kqfoiadbR1B69IRBWuJTSnFKZjl0znFFr
0CVtzIDput7iPU/6xfXaZUYyHYwL4bIJcs7AV3I++eWPIsNj5aWpG4U8/jHU+cEBj92OILJyMSBD
4Ew75FGMRDqKZ7A5qjFJyFSELQUcL/OQ51IqBq4Y/MD+bgk5CM1C+2eBlrU37nuKasKWS6wFd6u4
hXFivM+DKGjO0aZuE0+GnbbIamfUUzpQtHc10MdIiCHcqLWQr5PWRu3cPE0upw42D4VdXbI3wFDR
9Da9Uug9v93Z2MgaUEszLmng4yaZG/85hel3QQ3WGn4PY1IBrVypFP990RWn9qrPTMGRvJFoIA7v
FmAl3rMymaVe7sWan2E/T/c0YL4urpxjIzXyFg143syo7aRaY0cWVjUHDm3iPSlWLEOzGF7ciZz1
EJDBhslQWAGmL+hkaHz7dnsBFI3t35tpq18FBAfQc7EYLPI3/6ItFMHqmCUHSBXewrBJ8jNau0iB
mlPZJbS70uBUuSV+ZmswBqO1TxegnoYBy1dCPKN0ldOpnU+wrTxPawRoVDAUPnvxyKhTuxHcGt+3
P6zCtjci+WXrOCTnt9xpPe1Hn0wQl9TeWBCVLDrQmxTvaQkGBB9sy/Q/tDAfaMo1g6eO2qu6nbyK
MnSXl5EP3CjBG4zU/kmTJEFZMLzdlAy1NsFj4Ct6ReSbJ/+XJ7HA6l7yLjZeNhNQdwgzg3uPBAaV
wJj+J5XttBz3Rn7ihIUIt6evZFcS0LSkUgwyKh7y8svUMKRjMz4YtakSahqHChkmaIZF52Lx+bUW
SuMlYD4TPcMeLbs1C2nVwDI7qoer/29lZ03m+7CIf9fUdKsYu0qgKGvw4CC6PL6cUwGhjmsDX+C6
/BKljZdpCv1DWpi0ftveIvWJnYbNAXJmbNyXxo0zA9dZ3qHUEyLN5GUrF43Bpp6EdPCgRNxGvIfr
lI2BMsS5TddD1nx7I2gN4VhHXHDOOnghjDG2VN/O57Crg860RqXcli1MwZll23bGSFCDxDStZS16
1nLpwWaq6ex6eu8TpMZVnszMW6b793mVDHwwekIrRJIz3U2KiSjuddmwxOXYZ5wlseL1zKaDPh00
y62C4boc9f1w5fgA+lLQugwHClyT47/zf8ump9x6iPIN7h7OQyFBXW5Hf61/07vkYtoR2FpKaxsR
6HptAfJ+LWIUlgY3qLqzdzJWv5Q07GQTRi8FFllP+xYIeB+DV3MVa0HFt00PkegKnelIJRMM+gaM
HnBXrd1q1ps+H2OcdxCwarfnQovQyutdRJxED83KsZGF6H3IcgcOvVdEa3YrQHE+7ZvKpx/9hkGt
WlexByb2Rc7FSKolkIr65hW37zXLlUizfpTUS3jR8kTOUgYKkAOmSCtIecTVN80MhsYzFRHeTnZ/
Yte0VATSY8oxI0D5Oc0rG31TjcLXf5ngQnUPoX83U6bU399Op77dtB0nRjn5MwFkOXCtg2Ntyo/c
iZ0twUqNXC6XSIM/Un1j79GpFxNQzQWcpnMEgQwaEQQpqr3PpdHoqcihCF75ITc/p5aUrfq2BZGD
XkiVCAyYYMZhm31Rfie5ShHGFO4nIHJkfc5CIntTKB84o5EPFQY1iLLuo3QQ3QDWnaSEPVMq5SkN
mA2srnLX1+SsxpKKvOajIBFo+aHpgu+xw4Lp+dnVHNVqXVJN3G7k4B2fVqRlnp55kb7oVdtLOaMj
g/JrX78pkMctyVfC3ijt3Ak6QzDVAkyyHvYLhhzgeHy912FeWsyMs5SxJrZe9cLofJzkUEDURQwB
cIW1jLVxHI0yd+SMVrgUO6JW4ibBRwMqeG0Xp7Q1AiokQ0sZypOJiLYEv50yG3JBcYHHactzQwhO
wRzxCGW85hmP0hYFfVr3tGR4lV5ImGhncmkDmCutd6lOkmMaP3jSXUxW5bVnFrgxEvWueAzSvTYs
Lt+Q69LD7v6oue0NzlBl174ZZhU5nAoOia7MqcvxMe7FDgEOueQ8z2452k3ynakwt+9ONZaSLj6B
9ADOyENNQxE60jstFnYT4XbxYDKdpMdoN+Fu6px9ETdFlDErHSYHJirsjZjE6WhCTXpblXUyKOTv
+qlfywqbSuf2K0QK9giRfxAT6G6+fznHaMFv/J+9bfToip/MwDOkKYw5R7YhUZz3+LNghVMm1HwS
WS/iZq4aA25XEw8i7c9+pm5WonEYghwi+DWAMp8u9keZQpdnLlqSbFOpmAiywq+7xjpMVg8F+NKZ
1gdDFNpDje1qgiTEGMin+xFyynfCDDzlRYCIgcG+wGUtp5TF0KEDe8fBrmVW8tK8hYT7xiQF/H8B
l95w8YPgmzgSU0RgNZLn2hkqHJqa9Q+JPM7R5vmBGw1Sc/6palxyFBz8lJ46cbduYT67u/UIZgps
SZAZaiYNSEB8ygMgMoM3pc2gaHDK1//hYQq9PpQKu0rvzz96gS19xLhDMKJlbqxP09JbWWS5AOu5
qlEyLO1NVeQLp7gzk8p6HL7UsLT0uhyJNIVtIb2zPcvTcO3rlZN7D9ZSVboaJUEYx1GeXNLVrOI9
N4LBsQ8cB2Rm9FS29hDN6w3gZWPtgv9YABtPZeRzbRA9vdu+fKXRdCNSLEW4L87XXI9MOGtcXFcv
hU8GE7uPOv4wqPbTO40KWeJvrab3YW8FnAgDfuL483uxT1FikdvFS+QuJuQ7r+fuZYhtfR7YLnZW
IhHjDyzVx3Q0iS9cJA7EBwMiTO1MoXg7NJ9u2+L6+pGbZMlXQibwy9InjMQTuci5Yyu7zzI2i45P
LaTAzk8C/w4KNhh+WbY3hjgu1COGOL0vuqOdg3vR9AyNY/ZkYdq7mi8Mb9znju+K8b9hcsm7y65o
is64aHvSba6xCePRMO+c6Rf6k3i/vhrcAgJJwued8b4NJwFypZ7eLZmhPYPPC23cPWrSw/I8Bk/p
Cp3LnViNmY+wtUe21wTv6EGrcoH/1/RdadscexdQQFvGVB0VtyhaW38uUQeUMerrAX496itonkox
t+aRxI7NN1gnowAiiGo9P+dr6nuHobDoKrNF363LT4UEqVZCj52XI10QJmOPeVIjLJG66mq12b/1
9d9Lq9vzfRgklvRPZENlLVQ/zD1iI899niqftqhAqmpRCSju5uCStwPea26txgLHJ5NhVojfxl+2
9mFNDUwpertP+M5U97ydWbxeTvlK/AyjjAiq9pV8e9Bj9BdQEwsUS7lbS/HPLZTI+FHfZ9S1CXPR
4PD6O7SPENuuyR5nkDwx6BN6HocpoUw9u1+72jZ0CbNMOiHaYiRLkykUuCeB41WFIrE0sCt2fO3y
JW/fldoMy76g8TtZhk/5YnwDHfuIqdjHUPtGYZ6R/hqJkXjkLTNt0+QHM6gEhG60rdPR6WTJCPHB
oW7FY6JEW1SB7yItLHh5+aZotQBrXA4pFl966kic5GKzyI30QND7KbL0aCtvwqOZxI7r21Gn9Hwt
kP4x3q+UPSdoS4qz4SG/XWC5lnHW7TPCBgbwc/Ku7+ZPITl2rP8zzW/ZUKkfUBiEllB9EGL1nO3o
fMupuKgsncK8DXc17tU3FBwRc1kb8ZKYKS9nBWxPrIFdu29DMzHkiIImemj9PakQrrhh6+4XTnZW
1YIRrosmXxz2nYUz7O7234+TJ+x4wfw86vRf9rGeEjkWL8pWGkBWU/5qFwNAOfiMPqydfsbfPLIu
Vs0h4qqplZYJhzKJ34ZYdgvJf0dkm3nnhwNHVpZ1Id6iXbW0hWENslJ9taKhnAXl5BjWD4YeyFUC
Ue+fVUbsnMnybCL8hwBBUfCeMGh7MLmGBBLF4TrN6h7fJYzh1ryoj8k+d8OWn4jwkuRE0Aye8mXd
34HtXkOSNRwUjw7hLgkDBUTlVwlONdnPtJs+oET+vXtYVvviXm4VMlp+zj1zLT3k224RTABET0oN
xs84useQg0cHKB7EY7S6CYaNU9YrxYlPPWAvnPyKA4jMVbkSvBX8F7wGAdOfLJbNoc/XkH4llDgd
TRc0H+moqQ2/dHnxrQ6UzkGyKkvPjWl+gNi0RlmVKEnca9uYJHQ8KN2cjdSDOahykF4Y2at3O7fA
wYjQhfpZjEPKuHKnyJ2wGaaaFUXOZErQ/VQH+nSHFO5pUdWAswpZg/mpJ3epWKztFbyvcuRvSVnA
Bfbonj0D0ZoXhOhZ+sMO/tIQkVo2dlEUmNBujrxwymr5y+C5l6KhXJiMyckMT5E4CKiYeL9ZF7gl
OXWq+c2sS8An89HIxjhcNTN74S/SfCT+vigEud+zUVtSWS6J7NIQCLuIAXdOXXSHvYoEzDWbK1l8
Lu3wTFa2aqEOHWobDwasAbg76R7jVaii6yeXTzqxyI9q1Yq7BjVeZAH0gtibU+qibnK0/IL0a7as
uMOFaCZe5N2WfddeB8e4Zwzae3BqXZhDZlsNk4QEgLlFGUNHzhe4JSYLvYw9Ml2vWbEBDg3qHo+M
kM9C9SqFGItB4MT9W+PichJJ9zNmXpknop83LY5tka142nm7gmszdPVwWHzzTRTPsq/HznNFcuRN
AL3vZmQF1XwCBFO9KeN5ene9iiXVRZ/sI3YF5bTQSHYSOT5scnv0Bnh1KFsgTkbKXGucMJr7RTkg
AqzeMIwzUApUgcgERuyYHFSCFD026xcw0njxvRiaipIREuxG+oG3n9G+85mmbcUuIZ8tyWE/8ZyW
Zsog6thEVf1PhFQ79bIOy/ijhFt/swVm840vl5UF8MoS32Q9krSkwt8lq34RoKnIypLXDD3JiZsY
f3HA/+Z7PxooxpjjvIJZ4z44xvl6X0b47cuFs5RtPadfZ9F1TKUpJQhn5RS54kOfg8HnJ6eAnEND
qz172II1M/jRq8wa8A0X9Iaz2+8dM/jNfC2rCzvobwy/sYOkMfeq8T+4puL/42rKsXNzvDverBnk
g8OAejkFWcuuZdMD/pFe1fu00yMe/1NDPVmmOZSQtWGo9YNnFARPL6WfOXiDlg4zUlPJspBOQSyW
DYZWmyjIs403bSxlgDhcoN/G2s3jxz84S8K8w+CQQDPr1NaM+St3jYB627N+mvkp78Hx7KQc/o71
d7DW6qMpQRhq6v/+dZXWV5AKNnFGQZU6rSpCinnS1WqMyBjoTk8XSRNm8M6zYm0EJ4X+tUBGgC47
Jnhps/ROpIY1hgusiFd80U2XCu0Ck4IKbWcIEPqVBHEGrBiyKSKgPMMaglKOTphp3s9IOGC778oN
LeSbp5KSOlJarO0d63Z1jITLEj42lC4g/91mEo4coGtUu+xWB2IG9xbavQgv1iG+Lb+8h5JvRdXC
kGwa+bMq5rlGc+YxqK9hzCXrx4ORq1a3A7ayun3VbaCaInH+XTKaB0nWPuFsIJE2UxOMDKoev5ro
BGe/6CVPGh+fidTAH+RXFFOwSg8NzSw0zIjZFYp2cO+GiQAzjjgF0w2KKpuFsBIyW3tBZsWCF+/p
MQtIjjhIm983eklRE3OLFSWCFBZP3nIT44BWEGmt4Paq6Z+NuquBQ+DhtXFN6jRaK5Rz0u532k4O
sBBA8DQa4cQNKsk03/IBgr180E5KoCTYKy+1PY+WdV1JTfjMgHTwz1pY6JaNuMXhgQe8LkeaenM+
dtl+FZSgBw6f4IgKPI3+7Inr9tecl+56uKx+i0SUFKBXWUIjfpX0ta38ObrbnBD6tWWfyKTsy0zP
8tp8sq/nU3mmmylVjfnrn/9i9M13zbqAbDoDCemJrPvf9dkCvynxGwRlXl8XDAQ6+61wKskmTwcm
v0hYG6TbWFE7MM2KvyyeUPf7mLThgxyGUQYyNwk+3eW3+/uCN9y7ZXnxujQFD12549ECIDJzoVEH
pPkHuS/2ikmi5ENXXBg2uPH663v19X7eRTRuxZkxrbfweFT9XGxMRmS/mgtmzK8E00Gp8eCV+fCT
DT45AmHDThIzVSPilZNdnCZ0vMGrqy/dZ5n6dD6nsosNwvr8yf1nKYDNC5TpxFmK2B28F+N6eQu0
HOjZTSRJjCg0JlPHTZRLCJOBJVS5T3KE2YJAa9FYclMLNipPOqe1JoEWTfZy8gZf7GYe+m1DJkqJ
I+R0m/HPP1R9MqdcXgskKa8wyEnwX5SAfFzwu9XccKrVbZikFKJuzXgQp3bz1l1qVfKEmYaBqbTu
O0RfYu+s7frPLQr9zAbsBJKUMwtHeEMJLfpqgzSI1s4ieBSWecbwEL3/5StT1MtilSOzsaQ1DrOq
Ww/rHBwTt3SHucv03xOmueCthKA8yHlEQQpbcRGQT4fdNXEN+YRB1t4YybM28E9VLBclaP6pJPV7
uXVE5Xh12fs8pZaBBqYDOnoOXlDCWXM1qunutszQDrquyAKR1yDnxqMOtQBU99zrdH6C+t5QFVic
OqRswdBcMRYLI5qU9yEDN8yGXeAEIg3UzXv8g+EN2EmzDDaF1/yq5pAY778NwILhfRblf0rpFBEK
1AuI1msTJ597mlgvy6kiZFTrVyT/9qQ0/6s56hqDUBJYCNfD8PTqjXqNpbnwvh3TUQTI+RmB+jSg
1SSNl5ua8Fs8lR8uRXNrnKSEq/JkBbPHQj+9Lze01NUAqBW8r9qAOUPd6yqSBNi9YZOzFycWnpZL
2FQDl+3Ag8SyvQu875z5ZqWrnsqbmV8xkd5RJ0/HG+zJgYnx0B7IObFrT21/OXAoDW9NchCtNLZQ
vhJSaEe1J4nD1DHojskOotfI2cWM4qSsOMc/KF9cmV9aR860dKxsMHHIgVkOgTUORHegXRvaewFe
6pQfnl+Jodf/+zCgE90baDEcjv7g2LpEBoQibmbHck4eTT0Df85Z4GubhtC0jfACxHto2ez0ah2/
AyG/dW/54jNZnBQ/rwYulXWyXy+C9bO0kuXLke3i10JTKb5C263WBClmUPWhWLcF/BVnySYtmlE5
gHZtToppX2iaIX7UAfsAEGXGzDTbAePz4xu/1WmHLlttycWft9pLPZtYXd/FrezV+mYGWpsZPVO1
OInHMgWhedv7B0+JawLR2PEKciHDSP0bo4a+gIIZTyCDFt/rBsQFGrPsJGlL6d5zYSQb7d9E5NKS
p7blD385LZRbTQMkvFCXltswEC7fqbMD6aZZ/cBlLSn/J9E8V34A2gogfhjfyCpJJYzuzSuvR4+l
x4fWNfa4y+FGbQT0vCg0VZS0dFNBDc49mRyT2CH5T7vSVYLy7oVfXyMqeJSAwJkY3dTGuNLR4AFB
33JNvK2Xg2T2BawcVWF2yAW4S0/Bvdf7W+0MZ8UQspASWC+PfHEHH9maAdyinT60iYJZW5hlGpjP
OXs4ab92rTGnYt3sw5Vixj7vudCFjLFpnJmH0NQfZNXipm3qIABT2n3LgXbLqhPS58Le+wpZIkRd
FT3TP70amWbso8DJPhe0w9LA2hiCtWiLyiiUKll0HJvwjsRNxY/W63HY+cs8ehc0RTs/mXR2+LaE
dpdXkIzwWAZw7GpIKnhT5oVvnb97LX40SRSw3857Klj/aa0cWIUYWf7PwR/UUbSNc6kOBb7WfM/a
xsXPsbmokU/DcfifA6y22c+JKJEikEVutaNUITp3O+N1zPVoySgOPJ2P4ahiO24BuRoSthYngVAK
Cv6dxzAXfDg8QdD0MVBQHGfqj4sMXdgBGH+ni0VNmh0Dd1yfNdYIrEplhaFTxBqsZGnGBn/1Wp0R
DD7z+tWFzn/OlHDmCeBhY3U2WllKRyRll6MVq96oaQAiT+MMAFUEpL9pLRF4wf5oGvaQgUAqD9fd
jZrp68Vebz9EU8RV16iZ1BOUlmEPw0wa84Mhe/O7l6GKYiUGGaurOcwVF398nRi/xjjqJ9uec4p5
VJeDRHAYBfUzvr5v6qRwjPiyzqHLdLdpOx2uVB8xdWiuWGOmnl+XtEQZJM/WTRZGUGjud3iF5CxT
6zZSIOg9am30m4h1E/dECY7iZL48PCcXUQyiaGEf2HouADIt0JT9OxA0kptoBhhBUNxlM+nY98KN
m13VxgvdYZvz+xBfs9RrcrJJLrwi+QlC1WU3m/Dgh/ceFCekhKS7RDuVNCKTK6fpzc5WgIXzksTD
A9W2U3FWvHgL0gOgxhQdpPv1824xUANbb1wHcUFQ+AwkX2J8fi94X8Oa+eFqxIvHjDTFU6N2Wb2Q
aQquUtKDV9IK33DmgpySJjv5N9ypZ1OjncyRpJbvwrkrS8QkrNIWpHNcpBJhpzfa1M7X0Nqn4TrZ
wGV7+Jwnu/H1EpZKjd2UfxYbLoDaZLq0LMXodTM2fD75BvjZkPorRdn44h4s3a0yGt8TuZkrag/Q
fDVieOiBqP2kOJ0cafe0vMeScPn27AFDc4LJmspgeJxQ3Ji6wXOA/cUUEETDQyE/jb9apyt0PYeR
jb4BhDPHepRPN5JnWJil1Tr/dg6p4YFlsV7DxJsYsByaM9tOFfCUa8hT3Eon6Q9vEnfR/4mVWKOD
BZXYidMhx36d2fFHvKkmQ9eKe8sdkpz2cBwkvf0RkcMH1n7HRPNcG0phvUd4auQOZ820YC8DOwnA
n3jWeA7Y1cvnBtouUhqPM+GUGPU+svtL+yh/2FhQVIz+0K8ltS9vKqrOU9trlyD9zi60WlvfNHfx
Cc7Oi4DWza2D4FAslV6jktjF5eIFujAUgaR1/yMnONcAob1T3VEI/RAiNLh1srgs8Jdr9tZGvA0b
XDTwvmzgOWCBUKZ+fJuh68PMVv5PSNvVgiPmVnEIaDpX7eljQr+nVMqoRqCImFF6CNiE4w8RaJSf
a2BLBer7Xw2VkIlBOLDqZ35h9stuklImiP4Ak2lzlkkYy+wZqPy9zTtTeqvJDE0Elp4HCTca64i1
R9twXNx+fJmKlCsC1pk8M3QGOIv1Nf4UdQFN9f3i6QynezLrT6dbLVtShOPq8AamyVuLFFhoiI/h
lxS0/Ni68ceXzu3jric43bgmj8+kPjrIM2mVoMDCwnif8o2CPkq9XRowOw0OGSL+gKiH01XDNeN4
EBfXvkKvrt5UYOgs20LVB8yqn57XnNxi/ghxNue8P82gaiHXLPgMWxYDSfbsR+mfE01l0ctbB+Tx
i97o7+GjwNd5YuHQjESq37jzqvSIoML5p3LRnEOUHt7k3ndvd+zCWeJaLhpbJ2zAcj/hMsOUt9K+
RqDTBeFQdwykLIGV61yLv1wTZm67KOL1OIXMPZ3RKYhe3N5GkHNVAwro0ROR6C+3JhQ5Zz0XCDSB
4GwoeNlO9eUwep6flg2PFDcaYYLqF/8HfhKWIAq1W7Y0VQb7yqdj3uxWPUeemJd5lLpJs3ihBZiW
2/RXp3rI7C3sI7ss5/MSh58iGkj1oF1ZM3tQQQsbpnLMDuERWS9A7xfKq7mkHpFEyB9Me1Og8hHM
fSayM8U7Hs13irVpEPSq3e+2pWi42/P9LJb5HYu4bq06jszXsesML/dqZaxx2A7Gd+9LreE5gE3X
Nr4NPIZScDm7dktSPQyAlgKiU8sIqKvaOrsdRFIUP/Q2f+4FkrQYPo8K/ooLFxkPInkmiFb5D31g
MtbklFg15/Pdl315mkMWi9gR8i8gdaSrYUJndw69rk7+AGUTfGHvvWYgqJ8XpC7lyTwbA5emZmRg
MHfcFowh0bBVfDfeitnYzRDnDbRHs3XPs4dlnH8cvIZABt3yRCaVOJLhv7z5PN7Qj5+QKnJGi//x
h14Cc6bQIFhyYuCXudvzsLlAJ3iJur20fBnRceia5kAxAW5l98u0ioET/Ghbuz9U/kkqrRiBYTmK
XtXnnzNAk3u7Q8fm4XTxqqemueNIFtjZRLTJcVTt2kjJWDsFLCSH+QnaOTvavt8V9on6CywH/jAn
cC57T2mIoTYZMw5P8udl6NX9vDAe3M2e+jbpAcb0uzsT7JnciZLfX8AuzKV1c5etAUxWKMjPflLQ
32+osS9x30icrZasFl6C6pvtd6VQbphVNQJOONv3qEbSYUntp97J/Z8OX6zLCOZQQJX7QG0tHFQ7
3ArnvBWxNVixbrjSWcdn42GATStNbMCtgb+uGyDV7PPW2dKz7cq8KO81ObnpYyOPNo5gkbsttA5R
Clcnt0U0OxuAIECZkGEKMm872Xn3aTXhp9GJZ4iwKi/R7rFFwVNY2beiaMIHIqp8moDwcModug2T
cpJ39RJG2sB3dIXDhu/Q1Bo2pcBIsdAQ1EDVS4FAiUypzhhcfT6imJWlsU1CVSqsoaHcFHYlGQ3B
234e0fgppSAqcUfm4NDkhXe+5uSN9OMtgGBuBNgdBcI/nUPas2ohSwHve8T4/X2dGnGyPekfNhN8
LCdWUqBeqQnl2CzFn11YQCAXqEjBVkYHnZa3Y/JZHKT7AReVRkom/dYO6DcEGNGuMldvOOaqFUhr
c81fdJZh90aCXZ7mdllca4q6eaQUPQyNBB6mfR+p9n/kZDW2VQebDeo4kxKADa5Hic2HGGQzNgyJ
p2NTXobSQPRztcauvibWw1k/ogynGT+bBNDShgNzAO+XKEebUvU6ACkaO+6hZASGpkpPpN1/sk4A
xD9x4iVPbprCJOgB2O1fE4uVp/dymesTnjaHcRkWhctS4iYpbueGqg0vSGyFZ2w8MrxHl9MNlOmY
npDipfCxelm2IyK8H+LEIETM/uof2VRL696v08NuhibY8p3Xt1udAFfn4uxF+Do8YdPnxPP7lFJA
rpPpScz6KR/bKRpGtT1BlBC///SkLAVJL/0s+iuufuMl7wJ3AGKFUs8O6rV+QEhcaNXUhmcwtKFU
gIIi5AJTu6XYOFIg/qQGWQdvRPyhfmfqBcGXClh36SNegNXglP6CUl8noUDmRmtkUFZ4Npwyvujd
bUXILSP9rDS3ivE//vNTnhZiksJHplT+7Q4OLPChp5VhdNuIlppGthFbHxRPBlIoBl2+oupbSPpD
N50Wiw6zgpHHRv4KP/bCo8j/QCJhzy3tVSMfsRnUdeEW+pwNnTIu47x1yiY1UjOAOIC9ev0P6tjH
MNm9Gg+5D5vZUlC6VtwpQ74HKurhB/kqyehO25rjTxIINCT9V4gH4EEG7C0/qDt0OKu22xWHaa9/
QXhfigNY90BIUf/JJsyD3aG0dZoCn+Lgzh4wUiFYXqaIvO/A2/OiYH2nLo+c/wCVRuKbB00JRVpS
d8rUSyYqpCViWo9aH48nzctLeGP686qkLuGggT/dWjykCo2QAQ/U+9WhbbgdF7DW+m6QRISJl8jS
Viz+DYWTbxJy0HeA9KHcqWdPW65kNe47392+bmUIrKK1yA4la7F29KpDHcdAq9xtgY8tcyxHgxrR
JKpaYposIxdw1pS8fl44vlecTBwD56EGxgaVpVgXMyzQ4HDrzOYZLgPSImpq8t1Q/Quzlj/irJSD
3lgU4ssYKjYbFCDXGsLVYiAlqgqPusGeYBYJXpIFwkEWK4eMvw4RD1MH+d32K2ypFKS3ATfDvELv
lxQolC+0yNRDrfVBsJ9Uagsa3DP8RRnMk5RCsHOM2vMyMFLDuALfes/y/1Ks3OLdLs4R7dI+/EIP
heLAkTzAbnKPvjytSZZ41kfmrINM3OAaeEuLXhGx4g6XAx5eUnme8wcog6UnuZl2LIR/Il1MXiAx
2cVbYFDwcWok969lwQCbZ5wLWfhVgwRLEokt6tBGDCJF7peeieVzONgDy3s04xUy3MRPL+o/prCX
xeUEnOcfeyRKoXBgNMlDBYwFUixL+AE8RLsbl8vZunf3Vdju4hDDHnlujUdFccCt4/V8NJi/4PhF
Cgv5guzI1Tdq3YFW5B0V9L1LU+6icS6ZSUovZ1mcShubUNr07cQmUIOS0r8CGHBPJKFMSPaUHdTw
5fMwainki9wFUXrGmqa3tEXLMcL7lxID8EswFdNi7+Mn+tIqSSAO4dqwz5Zv0hIIPlq/Fi5CELaR
kLAk2JDBsl46AwVAqjSfc8lDw7if0Dc5di9OWh8pmG67vactvZa79LqYBHUmi/tKj0bhT35UKOxp
hEgvEQutnA0o8dto5xpLXQ9YeFXuIMt4Vinz9HDPIJIxF0zze96mifEw4xAlGDDsP0p5RbXIjnIw
ykWI3yk6pYelSSNSjLHnqTJYaBu2Ym0U6uEE+1JT5p0iqBivCkecmDHbElg0ut2qlTitMxMJtlq7
ZTM/y+xHmTsiG3UCtf2mKX3JbwPXQy89lWg/O6Bm+wkdrmZv7Zx06kZI8VvP33IBdRfLAOjsGvOk
fLZtynYrQYEMMvj6wTolJZ89Lu3O1RpTGQ+CaqAtiJm45iM0B2lRNu/EqdepW53V7zVghhfLuePh
Ajy1mlm2Vb+FhdkbaVP/M0FUqJlvdlnggri0KHV+tgzJWot7ZRaPNwzXtPLm3/4ox6+FgHV4jrmT
C1AvpG5mpz2PYvEF4YrdoSKjIL6Y1RO6YKJc9QeDMdLzTw9Dub4/stiN5V4M9VOk6ewe17Bq/fZf
SNswmsJbja2LBpKOHw1hNrt7irt3y+3u64gZPcGKzaK5cTW0UyY+Jay2EXvWeMcCP7csdjxPEBHh
Bd8MimAhbDKLcGomhoAKvSlOohb41ygE19pwYt7+SsGYIGlZkuKewZCynRVG/olLueDm3TTizjrv
Sj+HsU9WKt/3niYaSjE/PsjdOMoDIdzh3wvHJPTKfjlkgZJwPHwc+Fhm7yzPwBMF0Y1VP5uiSCte
7TDBby8aFHr2x5e68jC2H46tKngqojrORYlAbp1Bl48WbjJrtav10R0xZCdJyxXhWc9z/5hpeVFF
HYdPWejUKhUqjlq5cdF1wlKIvHwAi3T9QuK+CYt142dGxUaTF5rFezJF8enYuJ7oJzOk8LCyUFjf
b2ytKbF0t6HNtRxZIbb+TuzJIHPNe2AiAgFJCVXwlts41K6wmEPcPzNdNuQksTUhj3T9o9XW0Aic
s/lwTmOGkdzZ4vajYhM9pElZV1rg9OVuPQpHCE2NkDHg472y281ZKWbuccuSiUicH+tb3oux1D8n
3TLwkUl3EVC19hwPwW+gbpn9+Bv1xxQmjicp2nXXzX0nfjukW0PK2hJnsr57FBvpQt45PuJJzt4d
sWWtSfXijT01SgfHG5NTKlAMDYkl7VjYyVFGppU9tytgom931NdWdsgr7TrvxW3k/B0COVMEl3ls
n36EgmpjCju7Ckex5s7juV/v6LWWX3UUDk2out2M82d7bJhLfRDihJaI38Uxx23mxQnjuH6iAN31
PoC8P1eH0QD3DUrVgmxE8eFWAVQcviuDdqkY0GVuk6vGRafgYKleR3qOOTv9hfU+FwtCGRE2pzXP
qDvcrkRrpUj2p7oYjcszdh+SEHgasXdKt6wKkZSvCaaPOaNH3xWj/52McaXFZi5QkOO3ZAEZQfS4
Xx44YntCzHMZ+bUJQtJw/C4KyvKVIWmT5DlzDEnCLTCARPArbGYXBwzRVMMBf3WTWfpK+CGcuwZh
EVRR+qJ8Yz4CnWo/4MsZog5gbwQB+mlgSmYAPysge8I4Uolt5v1VlSYw7n9dOQNXb0FhDuh7ZBI4
9fDMzdbpZ3+hlWmKLuM0sXxiV5BAywGKtMfQV5MsvcD++Y4BvaMRbcrz2y6xJzHJxMlXIe9H1z1A
EfROJSJuYrMP4rZmWJhWolIhq1ryXE77P5oyt+05+/Yj76SGUwLCIYxq//tyY6UJFH73aXOLNt3p
oMjzLfysMcEggEpnlRwGQq/8V3P3MABe12vahIzBo+wbwFrYPhl1fNCdaZI6AyypEVRXEYWy9/ak
yocNSFMILU88gW7Z+cc6QfxWPle0YRbhsyn0VPOM5nKjo9SidfNpbF6lAjDlSrcHtH1S6/EBBXYg
CBwtHomft5VdoC8lEuLWqO7wNKT6/d1iU8d+oyQf+95qEZ/W1gJ2OYV51aWCj/FW/zq0PSF8HAm4
ifpDF4JMQ5KWZpl8iWJeZX6jIBe662MIu9Ehgn4YUVehuvPkHGJxA+dAWJabrIoizaqDMbi9xust
dTt8kv8r/pGIk/EMYziVntw4Bz37pbL//4VHTB7ZnkBugsmgjXbg3Gyt0oC5gFQSGE7EucMHSb27
Y9s1P/qn11WdvZJZp5FrBGAb0d5HY6n6fnnQiMerTfsY/35rNCp0jWEkF5VmE+KbU0sSVFC9T8wA
zqeTRM8l/z0sYTozdaBB4lCyoT/l53XNO0GcCVPwQ8igVDeQt+tGh/WvDXcuamBemHqgRSxF5qHp
bgf9zidEJTEfL8hwLz0DI9k9fhe5ECtGr2DCJcSRXskwPJ5+2rIzmC+8+XDuQzTpd1DhhhMT2raI
xtOn3i/DEz56RizgWM5UJKfgE6ISpXm3fMhH0X5WTj4jkTTTw7zuEX96tRfvOQRmpPetm8XCjv7E
MusftNH41qnhHuqCHaZdYTqgPoJSD1lw/9//nDX87iPUJa+oDGBGs55BulRnFVTSrZXmDKfZUubz
UJsztNYX/tMBhD+Qg2cw8xOJL8gdTza16fkbxK6MgftsJvtlFOP8BjtTBZvKRnQAPbDjYz9bYqJo
3WwULHBwOSXrqsGguWuyLHu/HwWU/xyM9Wl5XRrmAneNCKLJOm0RmOZL7PZxlTkb85UKATPPus44
KFofcv3eVjNu66h7iIbr+zDssBY7d5ewzpSVDZevinLL87DOhctHGoE588ba+Y8WTj/x6Fa8X+8Q
LYsdKFRJmxCfNS1adp4idXWFqyu44G4NTJnieWWGL/ltcDzKtF1nXe5R11RNLqHn/vH7RQrvCePu
SXjvHhmwwum4HZInYxcwyBUcDozh3IZz+kmyUYHedeNtIdBgSxuoLJmpOWLYRGSckHYOKvBtfmXe
mbp3KimvA4ZXpyl3hqaOhertTzMDr1eAVIMjyOAX2we9vysyexSmNDjcxVraf8wuwcAPpScNwI/T
kQdEzCxbP+3Q1AyrZj5ROIMGcmAtx/PAMsNNG8WKxUMOpxZZ/AJ9zWPtaunGeCbxbj6WNGPd3u5D
+9QsBQpCXXdFzEJEtSUgrLeinGKK52PUE1pDhW6iqpVHEycdT0p6RT0KyQPTqJFGpA+YuDZ8qQlm
Nkor5w7OzoaGaiReGDddCD4+4CISECauEh6DjWNVlA0Vc+TH/+aaK6ke2mtrLp34aIwvgxPaOWda
N//TnxYEPBVqIA2IB0rG71wa/kyBBvy2eEXg3AvNzxvBBelfJcUbeEhuyPNIZ50l+s+dwbxjc8d9
YoWLOYiU9i3ohmbAd8i39qftPxpnPUkgFTboQTOo9wsdcIRvSoV0GDtkwX+wK6AEQJAF0pDOJwGu
FJD3wx3HJrcYkT81I6G43fCuMXDSqTfh3i8WAFAQYNO4prz22LdJ3IMHopTPZCEdlYoSZ9vH+2Zn
ysnPoztfV26CGrI9ZM2vowHNEtybEOR1ZNldqrRu36XxmEDeJ5JZ1nHxlKmiIYcRlAlttFlaE4gq
APFMluQtNUEqA+rXVCJiuVXb1Alkp6tOV+4VPuz6eCxUQ4u/kQ30mxwck9cKryGgf5mPKkMtGCgf
HfllxgruCZ3HYJKASvbFt1tQhroX4+sjJ1gBHG5a5m5wLQfJnyn58PmVzA0l38+8+9g32MoO5bX6
/E6E83Jnb7DuTVW6KhFXVFzuOVq9dDNc5bIXGCW8a53GAXtGkdCbfcwjAAR7wrCWZkZwSt+r6rrC
Y4EYWjWi5KDe5aWkIMzqgDPy6nlb0NjtwuhbivH5nEyyqAiXXrL7VKE4brXV5M9Q+q387w70dP9j
5EEKNWbDV6P7+IbjIw+/stJJVrYvzKH0iUfr9Eg7IqbD8+PWCFQ7gw6sp2uCW37mhUaFBQgCCggS
shkzFd826np+GwWIoaxl64WBicKoZD5DzUKE+FJeHSe3P/eeTIjgfPpMN80dv47qI2VVF4aRnA/U
sHc7MxTnLv7I7q0oZZyOTjNA53IqLISABQw1fM8teYCgBrLh7a5Gkptq5NxHyoJ3OYeqPqQlCmcq
qn+n5nc9gJ2258D8sCOcJozzpTJakgkby0esHPffFVo9RFzaDApzEpLFsm5loOp0GzORAlyquNPW
LlIRGmAa+EXWvt0ZaoaQSxBJ3U6K6hziGYZ0ZiZ5HuFykUZb9rpHl/eTEfk4TbMxkUUHU2YBi7nB
gJzAtiK3hYmMuWyDNL4WhUgzBiX4ewCtmdeRMwWSr4GRYn4Wzk3AluG9yX+gRQWWuKJiSRorCKhO
SUUdvekcZYYqlm30X8iu+JHMY7bgduUbDVXnkq1F6HeoyW1Uvl1gsT6GTfjcfcSOTnU0M561RTuz
cyY0Z9c1eljeOiSmJbT2qMiZ3WAle3/2k3Eez37rE08VyOf8cQ/z9euAhE/JH5TQ2mQQ8chPht8J
MyAPPmsMNMLNq5lgA/giKus70fo2tfevflB3USW7BSbj74bFqlGYJN6C7VwfhL+nf+Kbt9cEXtWO
uZL5u0YAlMbhbyPb0J8TgQMqlgYUYW0ndKd6pRGoASYQ5SdiJeKFiQBYUsHJ7982fveIBnEFvB+k
KG/J3/L5h+++05ex9F/mYzx8+ls09pXQ1HNgxnbOt8ajNNba3B5vhGxvHIGDaw6Wnb4oWSRGq0kw
aEVAsaIZZBD0DRq4Ljq5Jcn0ZaeefenZy+/JQbReDU7vqyqbImzuNNeUPLx1kY9cmwvBPxnVRxyx
QWJM+C5ywoaZtcOfKbTB+TUiooRqbg/WlBj3wtJ1iXr9srV2OSuq1N5alLFEMMT1LYTnAyAyXWrR
7P7lx8AsF5+NOLy7aInCIfKU0kS7Ae2TO0xczXPdQjBQw2uf4yHd0KNpk36S0Q5h7KZ0t5i5ywrz
flw2WRr44dTeRSrA3R8qjUFO0lRL6VAh3FI+oA1Hqn+AkrD9IVFdcaZY1bzeQQbl6LOdSiczMIpw
p/pqNXzJIsQZK8eK8EnVbeOPcIwWGR02vvKMAUMbVk/BQd3WRknfocqr4slV/XCfIDPRSjjz8+9a
TZPTD9Ti50YfX4zPkUlxfv/UKbUoJ+BXJq4JmAYfFUiN74rSV8esSQLF7NaqxjJHD33AW6ZBOJ1+
zrKtqAwfMyWLxkgUQFX03mZigGNQkRyULdZofNEoPyzlp+d6SVGd4iomBf1dKMy9zoi6DkFYViNP
9lHvNIUg+VPoaWNmu4eZGWgkgc2DKMzwRbxcgKGlEljd59ZT/ksTc2W/oEXgwgtF7Zof3QUgrZh7
cJ2e4I+wsmS4frUHAcuWE6hwMwExv+s53N4gpoTjVJuADd4yFYMCAqs/DQGLZehCaOpKCcZn+p0o
2/DrVBlK3YZeJoK1ndC1woMZTow3C0wZ+C31xVyf4NsaN9JHdNPGMdx/u7lThznLu84KXaQ88ssg
/++VJ0AHXtyRenap2CMw7fxO1G9YO+8rFq+S3E3k1j35fnHGkt409ouF37XYM18thDmfE64HFDqk
yrdw6VZm3K8WjOgbDbE0TVw8DfVyK4XingJ4vzlQ39nSVS6sIateIb49LtfoGpUBm11N+BuuP6qv
1CqrW3hk51EJ1TkYFcG7MTUlxcZr0bJRbpZNELjnuk5RHQ5uw/1PUPIK3fLtPUKos7KWYh30JnbC
bgA8mFKoBo4NkuFNQ3STixmtnY/BWtqLdTY4i3OgdULXJTpHmLIGMuOT6rdqwOOAoguBJ7istXuv
cVIc1tMfGa284XK8NrRA9jpfqYynDvH11KNbliUJ4TAnk4fy3jvGhO8+2qlhnr1p0uoVSER8clCy
9MD+EzUfGmWMydCwZCWDLZaar9wmTUg1aoFoix6G6sMv5A5a9aI/85MkvoeDPKSVAfYowPvmJcbD
bXHFeDrCZhdl7lGMITSrB/cuMriNoJfchsrTPyZ9rc/wjQ6DiG6GAImWt0gT/eQtO/9KMzXxDKu2
Vzz2Hn1BWnP3Y7l+jb8GeNa4YQMu/H+Um0En8ZtQ0VeNcW+lKbhu0yfv0CSEnyntovQcuXtg5thg
VzJSG+u2WHmd0gEPqWX0sRa35sNuH8CaH90CP+JCUNbnMOTXwo+UEc8CC5BKRnaR5Y59AvrMLTAa
GiPirAYcqygr7GN6lhbMrHHVusWbjJHIZ53Nwq3rNM0oHrvW01ynMxPZhLwvKx0Z/SbnLvs35+/Z
CzXc9QfOHQvw1DHyCvOAufhxztavfYkUcw25KnlcbCklLUwIz9Peok6h/7u26+iLIm0PHg6fk1K2
TSYNRvLbpPxauLxHeMZZ7NrQpMcdcxZ6OTb6gmSAzhyu8oIjCUrsYGYAEZjDip0jT+fC6iqIHvr+
c47FHwbMVescWSSbcTdWfJADX0ottZnCCOmGe+8PQZRQLpEak2He4AKDmC+FHaxOW1Yj6P5iF/bY
ZWjSK0UIZ97e6GVGJ4CKE6TQF8bNTzHikYjhnQhTTk5swbFOFZxTP1A1O7epM1EgcDNeSNIMo7eu
ADzenFTh+fT4C8bs8O3sEzi/moZ2OELrqxf/mLTwKfBlaL/8+cjqgNbXpe5SE62J0MmU1XTzBg3r
ZkklB2Nt5bYx+PiPnXJD66OTfQYqkmyTM0csdh2W/Ovj3QqFKur2yC+NhrlMkLYvyHiyzy99tk8z
pLNlLBwq4fb44rPZ1Ak8VvAmzESLTmxGykmq/pESSz+V+vriT0ERfZE7WE1YsuAerzaz/tsm0rgg
csv4h8Wrnb0/Tl0cCflrxyVXAy4QaQ9Y/pKbmdkLGBpVVqixnvJ3p13/ZN/VUrbMXFvYxG5MnmHX
T+gsw0yWwZwmkezPWW6PRVhxPUrVUhBxI3oKGFQt8KKTQXcoG5ToiTGycKXp86kwhaBtGHaRz76x
c5F1fZiHxG6buwdFPVN5Uaw0VLvcduSIMZIXSs+wnH2XguEBhj1GWmDNpKj8OhElbaEmEPw/lhad
BjDJCNCO2jPZN1cWOg5ZEbDnRL3jQE6xbwt2KGTWbxFRMaWjnQc7LwKqkj+yQLRV4FPmSRd0BlwH
qM6qf/JCFUrTb7OcWP89Gd9+3R/kzaM6FYH0RtwCMvSQi7k1ANmRtoVUcwzvvB5GXVb3uevJPtpp
h0psXjd7S2IRyHWjIYUp0hJFmHgdQoeggUDmjA7sSvNbVVIfiSEyv+6jaOJZ3TiTUHXa6RV/fq3L
5+eifFL/K1Q5I7HeHIvBmgfKegjnCWRGDbXqN18qD7A+LxZoCWGJ1py3epjKKVKxsn73EDwR+vFA
d9cyiuGjzy0irm263uFSFaBtJ+24W8Nj3txK56e+USmRs4233ySwyZxGJEZNOA1yEvC4IZ6znmI4
CuIwSOGY2+plRRdvVOgw1w4WgKOoQFzFBYG0PFSsOFNORE45AOYUELKyeMs5kgF8KmxH+n/O19pa
pqN3Yci5u4o1hCHncKS6+DOa/YPyXGk1ZiBw11Oxfv9JJEAdPK4c7T6oZ9ZuXhI7f9Tv0naqqkR3
sYrpxdUk+2C+gZV5PpdEcTSIdwFSYwrtVKFvj2z0szljHODFUSCpKPJbCzv82MghU9CrV9tsLwRW
dfXX+zxckfih2WiMYXrS9K9dKvqLtHT961oklYS+iGvm+qRoLmjSxbxJ6gUteKvtwsDqH+4b34yk
jSSOs9XrdNZxOOvrHIaEMVXVbx8jXOb/1ubaEjyTrLd440cl886unA0p9bxY8ZpEglbHeMJSI+sd
Tr2nEICzC8BUwLiZkI51F5pXQSIbv2RfLyb4lzZCe/3ebB8M0IotMhbhGX+i2goQr31LgxNlx15+
DWTWksN2Sz9mJDNtt90LECjsiDP4nDy4xInE7H/nc2LLfvrTBHw9OL4fnvoOn9jjs7w+ZL7aRzht
YcBDn3xwV1MYJjsnM/pZZv9EdnpcZuqstrhzgfDTPJwHtOgjGHjnS7iwhitgTGNUTc4jwAgJAkbI
ofRr40bFO5CtfvzxxUPnYX/oTgK3kOAN2FFciK4Z4Fc4tjqnHu2S83b8RXE5/YzJBJcfu3jEktk7
yEnDv0ZzgA43Je3sIheBo9zqG4NRgEc74Uothdhfl2T/RvtCmrSk7yvqaajWnnIU7WbxL5uikMwd
WbvmcPrNclz0xSDuz9ckLgi74xNwa7HQzzrFSTpD+IzLWqXnFEFHTLYEg+mtFSJnwQ8Wx9ypdIYV
q0/wmEuDDR/VG1gCXENwhE5rviK9CX+2zq0dlbedoDtHsk9wMxqvbaYivbaaLLaiRCaYlVtJ85LN
HYqPSO50oVu4cHBQ6/50XaNKP+sJlg1A9+WheAImLVt1tM9E6mm72ECA+upW+eeIoNqcWuyB3zqy
kjFiDjlDg8H8Dht11WDp4HI5E3kAlxvL3cE3W1Nlmc8ivmF/3pays2qZqAadTk6f3bkI34b6GUGi
S+UGtKyunV5U5fOLEByczaZY9L1bVfx3fG34Fwo28lebHqL71SECAuWwTHCYoFokXHCTO8eX09lP
H9fzfMkNNKM9wzfP10v8WvFq4uqDnmvFAAvqNMjFaGiBjrka3oc2f6o+KB914QAKQN3zidx+i832
hgf4cGRTsud2SNhGXkEKbutkTkWD+FP8uoRiEiryKOzrDaPy+erxdSPCBR7EQjYBnSRN5D7ugNmf
RIB04FSDdzn3T38igUZ7TgVsgKUXfaDOSPjP6zH2PG5BlAlJ5L0q874k7ra0SgIzYlAF2gHTi71l
LSvxTY9Fg66LbRfGfmz5juJH8IAHgAgn5GQwY4JMTZdmMVOZjiJre+vttq8CRCDj43Af9yLblCC4
EMFS4cAep+NzvsIAXIVxGgv6/kBIre9lQASlX6ww1xO/OceuHLLx9Q3MJJQzDWDCi/9VCkYvIdEF
R2ugFuFDeGKlD+5AuwFUEylJk98d2sX1Ia3leK2IqmhV+v5wfOH2u2iXF2xbidCddi7yXsPSq8nW
Slo11Fhm4iwyqZnVWI8TgAKLKXlm5gZl8rjZsHJzgJwu8RWXoIE0VHHWtYL9ozKDoh/Sf81xWM9B
29Y4IeMV0vrJzs4EoSEGxhJBJlnlco6ZxtlE+crjLmCQ8liqE8WidmvtMGuZp8j81Bv8O+LCU5LA
LYd7Irt5nmDKu+khbaZq6M1iFxiUj6lcLFEyq6gMWkCHpR5IvCskmjtZP5mFPm1kVPCjTL8B4yN3
OfwU7bnn5nc+jqh+g5aHcRGdFuAnvl5NU9umYOVC3K2bKURWl4wT9drhjq7dHJBg7dY8mr+DcWIj
F7JP0kHmwiCryErAy1FS1SXcQb7jU7uIQpZ6A9ZeIblD7qo+hN6QDK0xMsG4pEoYrR/daqvvDpFi
JZg91y6zi3oNlvu5Z4LXbUyeABiY6axMlMdrpXiBKsTNaXC0E5f8mp//KtbboIf4O8k8bFasZjF2
/PD0JDWaHvLbBv+S/4wV5zTj5VpsSC6UsJ/JHkKkgarePCuq/du3BMVLNHbGPym4eOsxqaopmCTm
y2LTmLua6Wajtvc3Li+JYoYLQTp+L2m1XvNLTXKxTmTmG7dMVBzsy8ujylT5y2joHrjwWdCreSfD
CRSqUtMtAmd//ZSVNI4WqSKcV2jNliRt+/ut5I3A/t3QCbi+8HZ1ocYpjDzEsIRN5m+sLpbx6nX0
qbuWipoyA3kda6E1AyXXaLfqfzXehasvqLd7hl0K27b/9T+alfU/uTqNIsSLJxq1XSpangv/df6m
kFdRUD+FOTk9Sfr4NbWlgWpSN9Nm4TkxPhwcWOgrhXnZNfAzkR4M0/lsT1sHythswGfnWRe4b2aa
LIm0hteLN06n90xWksBX6JhTYavp4JZdN1wkh0LBJbj4TLGMIuJy0HV0+X/hgg+tlpwv469E/nlA
GNPz2Yhiw+T336e2zoJUyy9G3F6ckTy/vntNEZ64xY0z9JXCZi9/XfPoIfhI6XCaTShvH98YEvKY
gg6EANUh9YN1mU4s+rphCSeJRJheBlfIreJZ9I8INLzuM80Fo3C3MinY9aT/P5EsHCQDwtusYUhS
x5g3k9JjwO9bT917oViC6CvZgkQzhD1vNBc9m94Qpv1GfL8FkS8OkpJ90XYOpJooyqAfOSGOba84
KneqatbZss+JVo/nhMCCAqbYUo1ImAvK2pdRBIQhc3tpOd+F2+uc5mkMs1rM+RAQoEK/HfNU9SOO
8NZnpkq0X1Y9VPJnN3ho/SslGsa5h6nKokOQ2Cn4lPaEliCmpmi0lSsUO6jq2oroRMnXR/R7NjR0
Q6W9jeC1I3ItKVSeoTZ71HCmyOFBcBfJUaOfwgQv3SJsuKRFjDEqyS1gv9UNh2Xp3SiWqMtEVHKI
ocfCafcSHfxocFCVVH/Dqo4wlwJQTqtVhBp1EjgfK0Ovk1vkYiImDMJn2uDLpPAJDsGuqn5ehgjt
PRIrM/ROQmh+Rqeb0sa2DVE6fA3nCtqpuZ1ZJkdEFEiT7+6dZljxM8tw6G1QxJqSh6ScIFof7NYM
TVPl8Ei7TqHgM2n2G7xq+HpAvt++yQ6uwPTZYxjD8RXiRjDaoSes5TOJP65K88AqrpDpLSbtPSyn
QqHoIyGwaqPSKXzQHrpE8mPna3f9h+QsTBFRi0mfIiR7i0gQEvg9u61eiOLW6/bBTYf3mDcUZh7H
dl0HPSGIoC97jbPaLZvgV94t0ly+SMC7dYBmbK6Kqg9HB8PFOsOKcKLWHPWM8FnBGP1OQRelXF/3
RExZQkH3AIV3gjNuWkEAFu49aCh9DnEyt/RdUZ2ZI4lR5cAYAbVHV4g9Hd04d0LeZHu1aWOAG78C
ZdLvHcOFHQVrovdKi6FD8cWO/pt0mhF9lPC1yWuhF1Y5yQ+nvtjeIoyznvtA1QX8v7Nuh5MffyfQ
p3oUs7A4qHrfOiIsnwqnZ5CJZSkxV7RLUG8tsc6s94EyRlFaRhDe1OQRfGj3MMAgszjbexKZ6Bo1
M1mh/RHNcAj1+WvVAL7Lanfnn9C5npu5nTBTNbbKRc0dSIueWUM41yQLD14rqM8hOqZk/mKJMHqC
RH7DkG84lOZL29pRJlYKRgOvX8JYmEL9twGmowSb1jqWZFmnGe5TRAOitaUehZDOEfi3dAILzBVc
9ymxacEARSGQEPTi1HDISn2GUDv93sJgRit52sCzB3LhrltJRTceuygMwEpG2/X4sCYx34IliqL6
jRaTN2WK42z23GLnHGCKOjz8MYlbVaXd3RTD8v4QFlL+mtyk/YOUNWz/MlDO3cMtHyrjmkerCu7t
TFbwpiRRIBocjYL23RUVZ0EzPNIJ/2ctvOWNXh4+I5s1JFRlT94I8Wv5aLi4obXi271WFfGvE4js
o2dbjUgMXR3EvweORyHReLRmdKMvw/IdvgPxVkUHeXQEFThRPv9cYpBEfVrbAqrhMgEEq+w3PiHr
nI8EAGxY6cCvtaj6OfPv+ur5ZC4NOy+jHdcxClddmyG2eWbNICrQQZxEM/3qikVbmFJ4sDvIL/V3
PvIXeziIdj/CtpvRmtDi7Uipc8DuFljVTWH0YIR4I9PjU4jVm+GZm2S89cSco3QV5MMmJ/TnO6yY
aPX/O1GN9HZ3Jyns2JvS/9FOBlfK5bVmLlhnyFNx5NXAh7NbR/YYFf+8a7MSHlxqcGjg9zwIXY3M
vjbaQDP85RoN7KoAaSAsXjAYKV2MJhP//BF8krwj3Nn2ivuphvPjactrqeFh3xzF1B8eLe78HRbW
k8zXklf/ZFRQ5k4mbTqMSLO3mZKpXAfDuLfL3L68upLab5VRhdkxXLVRule9m9bzes12KUgPNGeS
dDmPvPHdNH8ndzJvib9vjyUuSjxHaN5hLWEXCnSKvld/UdqatbBpFoBl7Gepv1Tj+0VPZCwidI63
D56P2f5EYEFr0a/kq5Gc4uz7pEh1k1kJJzYvK4SABFHMcdTkZTKe5WusdCEMUEiKIjBxxtWYetzM
C/yDb52MDQGJp3NSx6JQpSBdAtu73NEulkEU6lV+fWLU5GZiu8civzO6TuU/ZocwBTyJODcqt0ZO
S6yqAggsObgtUWFjkSl6nAFtZVDuhrQDIlPYo82wTnx/y9Biq8v01E1Szwhy+C557/3xjiMZqUXP
7lgJJBaZUAl2/hkGnUEJG+spdJkI6UDbp/TQFqDcduLsluCLuXywckhhylFT1vpzKMk6vKcz+cXY
2B5LuGLekdUT6BOrcAC/lkcrcbB9Ohm832SVBCF+1dP9cGaEeGDiIFJVcdl15OyiRxXGzvKteNlZ
N+Av/auMbHiJWk2RH8kRuNis2OkRpR/dQsomaT5KyJxcdE/C3T48Abj9GU7ZwPNwkXAUVwVyuIjw
K2fwKERtbuG1zg2juVaYFnPC0DIi7BOZsZu4PmixP4h8zms2jiiV1r1z1/WKdHyvIfso7+qYXRZv
As9JIZiVUik4/8HIr+9aHONjkehjlf7DffXqkSRkoaHvOHfXhRIEe9rbMKwK33LYEOJIte2B4UqY
m36wUuseFrlwxkCjwTDWFJZQq1PQL7VaR+v4EAKntHlMxtJ+aa0+Ni/qSskKYvO316xS87qevstT
jeYOOz2j45xjsyZCgVHBljUAR5tBnkM9NNVbZXUtRShD5jszUfawb5z+eq8vI61asR3MUJ00wv2d
2H98i/oyvyK0LwrDKFlsbUTxGwkUVMEDtvRMOkoCU3iuPr7Fivbppngl59QW8dgeE9GEvLlQn6Ze
2ce737HMd/1fveqZBHVic5k3t0CAt6YJL2K1iONbxv4RpcPmI7FbD9XUsJp5R9IcYN0uYUOr7MUN
zPoHvYQm+tvg0HCKefnphC07h3WhUeSVYyQpjokiwgcQ/5eO6Ahm/k7SwyrJOarV2IKyULOCA/IS
J71LYToT0apVbP5yqq4ToVO7bhnhAa+V2K1jPFi0SIU/Y5XL/MsOgbyqp2vFjRSQyElQLxgRLhYi
z/q/4V0mK6e3WodmZGSHZq68HlnG6zF3etBOKwhP/tFNG8JdtLPk9P0C5HS0Q9zwko/+BnkSpvKy
q7qm2G/jVAZAm0HzoLsYhgtlKYJON5EDNtS1yDv/LE/S+yc41KNXItz5QjgOLXsGRgkXhB0EwRv1
6bkSkrTdaNQdTolQAN1qhv5aulFc3oWkjkTqqhLi/32xWi/myKNtFyQmm4p+jqTxdh9Q9d4uwRFe
ZMbp62zNAAfXR1Z50lY0FjGIO2w5UKLUgL6Y0eB5b7cQUCrN6ppOQMdZLFZqtSezn6pYpJTpFsTa
lA9rnnXOmWuJs1rj0VkkVnnqpi4+gtkuUfoIA+14ZxmMZP1feeH80W+FId1DIipP4mfqjg2nem5+
nORSwRbFecuRjP0LI1Yl/QXDeiitsbmmyl2RCG4pwrFuPWqigR5esRIxndngQ74CosHMWhhQGcqN
mEJEAhZJz2LX90WYu2ZJ3QcMYE9dbHoZ84TKtzUUDGzqbvxBZiaFBti/5lv0Vwcned1yTck0jnnp
e9WdQD1ZY7MrvZhxuhU1TfNzeRL1XqDpFewsTv1JnJCaCQf5GMNi1AGjOmRFglBYVeFfJej3mJrN
RGYUa3/hzHPEskMNX/7loHZ/aN4ZvVK8rIMYoiqg1k3a5uF66LxpVXJGTwtF//qu68qm2ccfAdAZ
w2VqWt6dSo0wm6yCAEbpp9jkIFV/nJnx3m8pKcRpAGuGQZJDPV6kXDA0/xZ0sh7u25wKUBWuze1B
hweF7zEdcUhshixrmwKEtW4FC+BxJx5m186TAw3ZVmvj9ZoahFtvT0K3p/m8IQ9aXeARty7eBomI
fVmrFAxOxZX6H07zwJR/kZub3poH4svvIxbhH7Rjqyxb+mI8DXrS9Kg0+RN5MuTUgsICsfZW48bq
yXdvLWFQnlW8bpOy+il89mn+uNszJpT1lLyoiYa1sORJEtHQ2oO2Vb/eg6IdznwmCZDpOHbNnlZp
C3AW7iFbEZLK3eNYJriMMjAkNK2vt5RWzv+mWpKdk7dvB/7jB3bbOEuYEuzXAXExRib1ih6hUjmQ
wGSvVX8EdvtNrvWUKDS5FXdUsvrz+UoTKDYmpu32sJo0ls1TooIqEz9VviVh3p8ceo15bMNGYyG6
TR2hKis5eMeoKmcGFqv3gZhMI2rYbuYbcmMeVaowh134J4BVDfjN09sT+arCt5eWbPLKt3z8SvzP
DatafbfN+cuKo7wzL7wPFsHQpSFPk61IQWqkX/MCBbfp9NgvibS6E5By6VUFTgevQ73uSbBwJLcu
CijPPLSYr+JfWah/X8OK2tatWiUgZPDhVPorSr/0FiBczP0H3QxxFJnb5cAtEITeQN+H9kmFWrCQ
yjLInBpklte6U3VQzBjV2b0rh4TlyniTOSQMWdH+RNg+bSG/2YwPNhd40zhh92HW83h9UPzGkbkk
aJWpyv9bWRRSgtAV3zcn/mCdPTUG2JfomkCIfZ6lWPJFVzjqdBrjuXZLm1iA+O9wHfUr65/DNmwm
tH4TZ1aCLQMkKyI9B1eCwHLm/mt4s9ZNcHk7N3b0pXlSc5xLFo0EvPCWGvS3Cybivv0mUb4q379Z
WvegQ8znjrP1QBBpw3CdSzqgp1AkB2gdEiBeD4lilhK6QYvX5/hnUTV7BpygrQ52KN2BWzQzWMy2
wj4O9M8fk5A5tA7rL6nonxdBmiYiKNNUvfBbAPEZONHe66uXi3OEn+RNqAs1/0L9Bkw57+GwZHDx
Os543nbE4B6mcvE1zy+EzSwf0LPbNjrWChpF8999cDDoZIPZG26WIw+zWeJH4pb023d7C3oT4IKy
wOYm42gOordEWjV7AtH2gTL1cYfft0thYFgUGYhvVFbfhIj3l8kSsD7N5XdaHdHLDwXDJ6/QNUVY
xAgm1P3rx/g/Zb3jTCUJvXnS79J9G4neOWmMRFJZ5rEN8pOZAigPiy0e6y9eV10259jBZ324lf1M
/wqQ/Clpl3N1wz+vOgdN4GxRWWO4z80AcM1965uOY0MXXA9RARdtmES3zuYME/BwsQi21LJddMuC
NzaJpWV05OY5+Sjt9LV280QZVySzuk25fc0bIaYj1ns32iwAqEC7D3vrw8Rzcrq/fVmj0XsDj3OS
tV+r0+ltZWu6e/BipDti7Gg4bbyuZcqyQI+In7nMKoP+W8mtZSk7s0mAAlrZ5W1PFyhcgMoOJq0F
+RI61IQiqrC4PO9wN3kE30eQ92f8cl8xBDHaHJA1C5QD33ScUvyIFhqppTQhR3fr+u8KUYSEKgHF
Tbx/NJm0dbmu/66g4bqnsoKbXoG02n3VmBuogxc+fL9D6EIggbk9arG+YzGxtCYv5p23suaZQiR/
2uNPOU/TV29cTby9nEBtujFuRlEIzfFp9+zD9U2eWkZuVEeXuwGhajbjlhKWcq3Z2dpkK/0/cKEl
FHJvt3AilVLi+PEm3QZZ6dIByC1f280eXYXBoEYNbd0to8UFbae6VCX2jNh5GtGqA/VfJXnjKRoP
ZTX8+C2yOj3fcP/LG6vh8HQoJaSsEzT6sVupl11UJHPi+C1hz8EULVrWHAz3vOFZvNI2bca/B1hr
bGuPLWG0rkayHPvenngtgU7/zwheipqosuFWd90zPcZF31cc5st9jTCnvVHfqrmzXVOyjuNIlpLB
+aF9yI+gG97mo+mvSKAAt2cpiGPr3mPFlHX25xADl0oJl0sVnv0uVlaADT/wjehsobLrLjbW4bgD
8X5WJ7FBIK6RPYOsuZTyC45iCOrPdcin35scAIo/wUrGl2yquRzePTUfsHg4IYY3uIgyBTYyBioI
RJ85gh3Cm0L24YiGJIiDWdFwJ7YrDy/fqOUajzfM19fFpQfwkkwQryDtvzhsssGzgb2Vy+NK3Zk0
PGW539NzEmt+/BDwB5+dC6VVk/n0e82QOlDmW+hREvkX99a6WyN01YjByLUYzb5NlT32Vi0efY52
bYmdfXIN4KvHuMiKTrkJB7esW6t6PSxSCh3eCOR2zt+MR965bTFsjTfet6B/r5BFLKwOjFyTkFqI
hhQ4nzlu1iSJ7TBgRsAn1O4bYwcNq4QlM3bPHfLQcolCMH/2tDYxZmxsXfkjMl2/omIzKFcLbJo3
McNm5iNlnyNRnJUZmH0MyAAOYjQtn7sAinDoPmAflZX4UUrsobdXCcr1LU6NV5jEaut4qoctj0Yu
2KSxi5L4ODjCR/wIvxRtHj3l6AiGmOP1AgKr2Vi0SdMzejZXa5f0MuDOEJDmdlGrN80ZrXjyWy2C
QCERqMr1pGifjfiOg8fJsuBLtIv/+iP7PIMLavLcCOKwU5YwrQmBTMoR5wca4dpv/j5gtbkK1ukp
kYXJNoS8CA5aKT32aDjPQRg20floppTOWgXML+DPjILM9Ev9Fa9WTs673xIkgPcDzudB4OcdSF2L
YFViYn923S5I7HJxt7ltx8kM9fiKCKDmyBqk4jwr2DNsibRhE1bPb7l9bavt5Nx+d8RpNqJu8CWl
fLInAS/RIjOaJzTKCGPofmISlrJAYFgc9UzDmoAgzTbpYq3xTB4trRLLhiG4LFnp6W+rjzMOTNDK
PYGAGffMXYnADP9YVDXBeN3yHtsxTW055JBOzHohZxZZVIHa+l9r6aEs34hkszGHnjVtPEKe/YSE
d4toVfXmdLgetw+VFHNrCM9XZ8kps2cUQQ5lWeaMp0Hm6RDjjy8nagZpPRXuqzCbQFEyiICPTtHP
dtuh0SEE2hSgCsMA3r2CDgbvxQq294OH59j+zdbzhhkKDvhpX/CqxuAPf3uUXjcHJY9f51NqEOPP
FmNDvCbcaYEheHjiFaj9kNjIamx4mLFWxBXJEW+CiysmMVO1WkV7pNluoDmjLMNTDwGtUsONr3x7
1glcZcGAuIXNGwwywNw+x6WAryt+oc2bVtfpqRwV3mSkkHw+0qIJJtg/N9Y+jiykTPsH1qEPGzhh
ZFculBG3z0+QsZHGrMOIWwtCaXRsQlypCFMu6EQE4YND/VTFrGINCWUqBpRny66VisVD6ZNRYQma
cjnFf0yj7E4oSxBP2Gcy0Pnac78FCjiKW0ruNXZK8cL7CBbxlkxhav2E762lhLMQAoalKGKugOTD
5JYa+0LmXVPx3v5lmdMbNEivphgZx14ZPqC3r/HnUY0uYz8sLc5uoCW2igUUKpEiczFkvwi50SYx
lkbCH+QHoAPIuC6+6vW+hbmvWrWc/q5yoiT6vgBnkWCfPmqWXkfl6bhpP/j1rzsKjXKBCifIv3x0
z3AI/C2Zx9BR843mIxBpBMJ4tqir2H2kxW3Bb2LNKE2ykLcBacPQOrX6+gJzv1ooXp5bgrGbDu3e
vMSVUZHGds0/tbJtsJQlmlNUXKHW5W+a86D+XxMSQCfwhj5Sr5E6lKVByjfoETIbvOYvtY7r49k+
wU4er3UZY6DEWbVWJoEdVgiEKQqh96NH8f5iGbbvSEmrAuvIsOCAsMdadaFgws3hB+U5c2WleCwr
iHWdQQszZJvN1Vz3PmRqx+U8xbfQMsHFmqzXy/pqac09dCanpo+BAmWwH8LNdtrxfGMBXVy+4GOL
LoNIBJ+Ut0NLXllGj4k7uhRe9KU3wiRYGAK3hr3UhKxA9GgBmTPJhP+wVxTBO2/QpA7A6jJ3rnAm
cMolgH2Sd601y1MziJ0d0fVjCptaKLQUPTtERZwXeAkpU5tg0lUdwXLN3aM7bNIzxbKqdSvihrwm
QcJFltRXPkAdyJizxWebLSfhsukDTomcc2/S8sdCJhw7WgvZTEIE4K0vY8FW38HIpjK1mfgYmFPd
xL/sWciCMvfdJyYYYnJqy4tLHoBoouwL411KFCszJHom0EFEv0LF33lpoO88Mh0tNY/xbEuxNh3/
//jyQAZMpUdvqUrbSEjOt77ozXX5SfYMnJittrmrSFPJEh3Z+qXhqU6YFld1lD7UYHQEvrNJNF2W
EG0InxDcOAsJD0HuHLor/bHWS+izU8t5ccyR4KYWz6gv2NJP4K1fHKXLSCPSDWM4oPoG3dNpwjGU
v/qtyVGFKIGL8EM+GHdLi8kP1kPJ7/uyHlu536rANaIMqP+h++7dybcwq3qDAbkhmeuF062VryKC
bhTnWR2a8zskiWIBh60zH8nuCJ6H6NqQaFQF7+n12ZW7f8Fa/Rml2hHj8kLy5fmHKO9X0t5rrsRc
09eN8SScxifFVQ3DUKoq0AZ0ejd5kq6hmhXnl9EACYq4vXpPWDdxWOWNgqc+cw6kPl//n4bTkYib
DjkdQeULMci/3kYkMKLY8njAOXUuXQmUeCVaG/2HWY2JU1D6eWJLPg7AKMh4VtyGYFPykM7O+jt+
0Yd6QIZ8ttEPILCA+Tdu62bZFiC+s8tvSADA8J/EGPwctZNgKq9zy/LCbT9oG1vH/syHNrMoAtcT
aN1zuTB6UuNcsyEfhxZBk3RiNW6nsuHlwBNF/1nB3etSUAeHW6sQu1W9AF59X40b5gdfpj8I/3AX
gYraash4/bAnY/Vfj1fH6pTY1lSm8Yx0Fl1628QR9NfK4kcNBFvfh67pT5ZPyNXA9pkdSzAQpA35
zxBDIuVsJ6tLpreEeZT0i+5Xicm0Sf/px4bVyWAadSnHbpG3g5rn8XCYHhhy4JYmhj5t8XdCpC68
2bSCJdYNIvSeRPaP0xnKqnTy7nRakphQLtVFd8WSF/72Jpb3ZNTdcwa3X9E/M7ll8seROOsO0lGF
Vj6+4hv+fggi23y6VwsrQyKUka1zH5mYN3IgicQgDMuokzezcYK2QxhEdLUp0zVZCL04pe6/m6pb
RbOq2cQNlKWVZgDD+gHw3Sj00xXnkyw8y117tSOylfPRhsLJHRsUCmyPsZAHZTZZ3lxjigl4xq+w
lnKdsLng4sOsI1K+Kmwr+WZOVcZ7+MrSxvv3VexDU+jfjH7jCw8xLxk36+c8JTzMcb1wTWEK6gRA
IaZ8gl7XlXda6tbIFWdKaqnJxFnxbqte4pzQozg2eeCv3UI8Y9lFVMZ8B1Bt8dSPusya6vZA2sAW
XgMfHMUmF/t4QCS4VA6xz7G31vz6feRmHzfUYB0+ppbtLsePoknC+qhbccDia4NCmcxSYz9HpWfQ
7kNqr+Lw1ZbWNVb/Ttu7A4aSkORAE76mtqQ4uxsHU3cbA4NeAxZ3xWVgFfAmmd3VJ44dhDx8kKre
hLd/KYufZyRSBmhiHz8I+FoM9vGIUbgB0DBDa0it2bbNF2dhRQbf300MRt7evsrV3C7whEDL3ldn
BmYr2DqFTGd3U7lHIrRGe85uBUdh0mc/lrFDuzSNjRG3uBdb7XM2uGo76c1MK8i7YDTYiY09QBKy
pwiJtKs+ZryqEX0nFnSkKMVeOpSW3BslH99k5aodMEKOa9fZC6LbYORe9EGgUBkQyJj0al6vtaCW
/weILlxastjWPE+8D5gP5JM3tVGY1/Gkfft6AlNQaZT0oGqGVn0pQuHRDfV+c02malSb839JhjtG
57HGd/wyWqq22NcmISEuB7MysYpVAifCO8SduBI8S8igo+9EczVHOIrctDdAYvHWQQP6djP1r7XI
0P0t/93IdhzJcRE/6+VtgxKHaIfqFBuMsHcx0LBRpv+EUQFSOxA4r02r2rbxK0GNBkpnjkhCBFvU
HqKrCs51aqcr5LsIJAs2hX275LzEPguDEXv5UGajKVJMZotYCLWutlgqYfwRvKK1i7tdg4j4z98h
7oleSf4Qj/ymleVrfku2qxPPwx2/+8lVriD9LSsX7exlISImqCDWMCqrPh0bxlnLAmRANRVUcmQR
IndEwwz4EPshAaAnGpRCzBnZYy6qRSpetjggr5MFoDqmQLmWdsC0cLqe4nWcwVEJSv21iTr2UEpm
dv7IjkT7avU0L+1Oqm0LFEy6g+ClV4zoJIvxArORbqVnB59Hv/zVtaRg+/wu1J49ICBYtdPr/MOj
MJLCU8/jWWufKoOC01T0k/DFuFIbqv60Aqj8av641cgK2UnK+j+bTy/ajNm9C1CejZw9JoiPTEUD
xzl/BVrUdNbKMMM+9ket6saFO5ZJuHtB46omtOr7zTf20Y8bMnylY5YOqXDmKH8JERCIrkDNrWeF
b+sXEdzxld4oI2XTNv2+5xrZkilguxwVGKU8x+KpZGJpf8NEx+3zvUku/aXODtpxSnW1X4qZ+8Cb
uwCeQLpGRGY0njwPpgY+wS5tUrm6WgoTzZ7hY/Ecf9bxB5yEQO062l1yW+K8lPx81t3eDgTnA5FE
UpkUyBNU1HnBi29EyetGSmUhVsX0AslfP249N2TXDzB0LOYUDR699Nk7mDrCZQDqYb0fYjDpGlMl
W/8Rdwf5LLjoIaaRJ+GhxSXSw+k2efGiErxi9aHv4uoopCXRCfG1k6sAGXf790Ixa2Jvgg3Kl+98
ReZf2A9I2gfQbafvPXnj1KUoQsb3fC6qQx3wfEGPT+fyEXb+DmbbOPI1goYDyIIq8sJem/KgOcn5
PwyBVp234fCd9NcO4asqff0k9F4cmeVABFkxOIVmyokjtjlHURJFtjcO/f1L/9Pj65qQJd5yEpej
AwfS7seMMX9+rQmO6bNIhnR1rzGOawJ23i3TPqd16/5loKvzlLRxiPcC7bxFMIVbRjtJ+eTYmgCZ
QBFoR8wzFBIie4IOl/jTJBSIc7MjyKbOo23z1isM9CNlbUyHqX/u/u4Pi3gKeC/89AV64ks3isN4
czjHHxtmeM2WHOZ2fWNHtV2b/vv1f9Wp2GX0m1grkmNxSy3tlbdt2YaJf9JkqVzavpnst/h+OBnb
GubqrcYkrckC66vS4wxU1YrwpBf1MIIp4iP8mzY8OfK49cfJs0mdXYV09w+lfO3lRkrGWCxqmCob
zjxxOcl3Uxdt0R/SXLQvxw5+DqFU3XD0imBFsbMh8zFFtYRHT57weRvggO4tcfRlVrSURfl+2/4T
S4YlAEYXY1Pzq01ChswPUCABJ9sKUDKgW7GN9N4fFYUtR/HxvT6c1+KUus2QHkTepFGWON0tdFHp
XjX1woACEFDpDykOuq5oHc+hy8JUUJddcuRGb13UqsKMU9ZV063OHHxymNhULf1RCY0tv469AqHW
FQL4Bb9natmvTxYoJxDm33HvSYZ5KhrTnA5EHctB+sCJZw70MPiS8m2lTbtjs5M9MiLv/OqzrVI0
Cx3YHt9+4UQO70TiYeUKqNizHJUjZNCyqdUj+sqyuHqqYUYJgefjNqytnhr+6nyuiBiEyf+NpsPK
iOlb5PJ78qrKwODpe79Oiu/ODCHlTHjKCCBOfLNgS+VdiB9u2xV2/PAsO23xIokDa/jOFG0Jgz0/
J6mw5/lZZ+QixvWEcTf/2JdejFdPKkMNr5ESSvgM3uBt2yLDei7hD+trVbwNUKXBSG0gEDv73iq3
bAymut29w2yshsMveAa1wv0OULXXw1zrzSJ7aeqyN5As7aRoVP9qUTkDtjndo2F4fzqp6LGr0fU4
Z0Tw+81HIDJbYadKXRQuHLeHTjuRbnFgv6hGCmC+U9/8M0iMGi/N93gggwjmiQlbJOEdVUfP1ID/
Pk+heSpAN5CB0NYwz7siewDc8uhrslEraK9LrrBfqNZOPyubCgv0XwFU/PrhqPK/PZx7GASRcjcb
sriLKwGhi7mx6j5TzNUSiFxFZc+cATojZ4V8iK++rCMfVmiT2o4ybQDsKkTCF8o6ShieoyjPaow7
VuxI+9FkYjWHl1z+0g0wfarwcrKA5tcA7DflNW1XF+phnNODiG4eUMhxTlc0H7w9RNeB7KqHNouu
zpWMQFmnXnGYKdZtl+lZ6GdLoL9kYxlV9eK3Zimdtd5gg0TBwDiyPENiUFhwLdgI4sqkZtXXwm8h
0XcZ2eyhCSmrpNJilHDJo1n7yEeuVPJv0dMirqj5qBMICWyBarcXpAJTWHqgTphczDaB0VNQrLmA
iES5N9ossqOqbQxbfcXZ66L5gZxJ9PmZ+/MIDtTVe8aY8cFpRcFLM1VjcWPGSKeSeUsVOir5T6TV
ddalv4VGMA8hnR9j5bxM0kEq9L8dVMd4HEgHxTBQWO4R6BrfWgNqKDHiQJiKOu6TBbeON/6Lf2/P
AYjEQmtKitZqN5w4daNq5Jy8wMw433wYOwTCv5I1KeT0KoqvmBQ+zyagzYx2L2czjXCvfRosrWFq
+jpKoNRW14uth/bnSt+UTrHAhuUQkFTKLdNfS+GwAEiruk1HbCgnEI1rPoI92cIXbOhA8GBmYv2M
GlEkcXMTWehRarVQni7Y5QQpJR2Pc1qkWViiiNgzsNc9LmwDjKiCh9YlX+3C4B8SmVhr7OZQWg7D
sfVot1e5xidizeWwXZ1SIdfYDkXZsoblTOYp5K/kbgYEb3XwPCKaxMvqVPJBx5Wk5gTV6iSUqXHL
xce9f6oSvIDsjWqZ0JAS5g5ac4yLTSwGsXUtRARH5efMHFIP9PDSQSEJWBAQcX4TLxpS0HsHQD0w
KBISedhJ2bR2w1jqvvr7xjqFynC3/HnLSyJxxqyIrt4MBODslFufqHURc0GS08ZhLfN09pVp03q0
6I4lcOLvPXJ8ZxNrMLJ/huIeinxy0l+BFSPwtDn4+EYmCzK1UuPiLerfd65FPrlrAZwSjlitEorU
BPa3pJUX/xPNtQidwXA/l0pupewctds5Pkugs1Q5jyLFm+Be8VKdL11CxTiFpuuBtY7/giKa0049
+eJqeualyv57a3ZZxxoT9j1GvqSNxMj1mfUSARHzwKu16O68kIxpXqcXtfpj7SbfbRj6MqE4wo1e
edfZQrV7PBmNFjr0N1TcvIUY+hgmZrndNHX8k07DybmlcBCUOo/2E+vHyP/0I+SWg9Y2oCBInzOr
UQLVT2JMwtaHbYjrRGhJ1ZgrkmD1SKOQXCEby2c4vy8N7AJjFLxCPk09UK40QrbwDZfbisttKQh2
ATvU6kKwa7gUkfwjYux7WntWvW3A0MmlE46o5BLLh9cqHHX2AUeKOGm7FwqJRvbL2QFcYKsGztcl
qDgx0T/EVcvjmxpsqmFwDQHIiSBSNIWdZ/ijn8nlmIwE9djRMbLFbe8sRzDIyiiF8b9H2atF8i18
Nv9uEM2hZcVH8m5bMK9QMiRhtE+Hh/G6lOGDTXkhgbv52VHQ6ns98XNxlTnqMIxUdtEqGr6/nLYy
qlIX3rK3R1Znxmx2+/QZKGWOSXYlfBH2SxDGEOw0eYCuq8sn0JCEbLjBY55ZWcfyi58etU/zeSlY
QUJQkKct+4F+dO6N3bj9NjiLveuaq1chjnC5UKdoLpDZoiXwIX4zOCxYRNb92CtPbR1bjm97mZBX
GnKFVWp67dtJeqIwN6LK5S8n+MeYipXWVlQWYkjiZtWGuFb1m+XkK+OIXXXvG5C41UHNJHcZs+QO
Y4A2axTvIuGD2MNtBYx2LWeW5HCCHotmgJZJJUWTSZOqv3aJx04/CnTwvcFbKZfuKsQ9nNRRnZla
D4ipviM0tFpgeqfNYg7O7y/0iXUNdTqDQ6zn8tCBJ5xyG9/Hl2zSrJ+8rYiRmFV6uIrL8ENX3vmd
LiUO6GOEiqsdVlSSnA510Spaje0SGmllLgezBbhClnklOjtSV1S9cgXGIsytOYyGxlI7dfqaO2j/
gFiH6nv2y8rHOxFIFuvoijiZk4spd6NaQjpS9ib2s8EX911130EXY47PjzRiEv6bXaqlHbhFmLcX
AmjuuTRQJBtWV89LiJVeIeqVNC8qDgLydYyHMPx429tAzJv7O2OUvzAJBMQ/51OaE/UEXWXchCtR
tFeumXAf8BzbqoTKDVljdeUpujcqqeK7p75WfUpIDb3gZjAFbbWcoPobR/MiLSg+xQJcwNASg7gt
yZI243aqIvTVhX5bo82psQYpQMncKnSTNsQmBbYKUTnELIyzwoBJppdTGOZvfjazkLmO/9fsmTsl
xDxyUZeJBlzmq6QKUdsZmECv4t5hNjn6IfTJdIBw+IkOqTIoLnG/bktSZ+S/4gAv9RE73X4BUibM
CCUP+lEURgKWC8yDhTaBg4j2bSMOhbGnc91mjra7iPdrKODUprczN02qY+gYZjN52WlqPf6V70iB
UnJYhRdU2E3He88J9GYy8s+cvHhO6peMYguAeQzqScbIvOY1DukWIGG3R/PMEA4xuy8woXZpEV3S
M8zKylTmRusQcLCnatuWzJ6DbS+kQQTYTuGuL5ziAIgTpSQlRdcZwNTmH/pVCytqsTNCTCU30l9v
uPtHyecV9T7OMG1rtWsUXmHrddR6y8fLMoTKiFD0SNduz/6FA2lvHAODWOJbk920fD8yyfqop+8g
WcGG8zeMz0Jsvu0mm1z7IcAx/dgjRL4uk5t5PfFtIdgNkaNRSSks2zFwdxDYVhPOZBoAn8C39oQf
CEjoiKjWszBG7TRX+AOMpkLOuRSI/sYrKMUMd6uFnwtAS3eulmRkUqDud4f4N8HRqVhSEJgW/rXc
U2vWm3HaTGfd9amIHU25iKWncSWglq5pW8sjJxnPc0Obw/GFMtoodUcoktgg6dXFCFofj8E4zgiI
ufXLDGLdKXTWDKymJE6TXXrfIlCchI5EMkuW8A0OpzKnm6mzRwq9trD3fxtl8MHdHx1x/b0Y8Ska
eEAkcBmNUPStCQ4CVYCg39ozNDgA2Pm+s8CYpER/VsVjvdZMAzx2H1bMFtdNw3w0+d3PRl38QQTt
YTu6PrVS4O/6felJySCcCcQTshAuoGZJIUKaKJUJ1EcnObn48WzDkm7KmCuIJNNmwqov1GNVJW/0
pyj9tlXm0JrFjZLkkbtLUcrJ6kOQ3O35qnGgQtaVX58pINtoBcwVoSpo+P71kUs1n5dxOdP9FuAo
wHqmvmCVSgsFk/aGmPXUhHAIVzDfKXcTb0HgE+PDIBVXqFmMekwVGL4bnjYvZmK+wJb28nrobeZI
zSVoz84bs5q3cSIUfF/JttaH6I0Tp4zIeJvhH8xLw9zuX09Q0llNWsepDfOtOMny79No7Q3pbtBK
g/Mm6JtsqdZjnXtjT0HiN1iTDijKbs/GTi5Y6XA3AudXuOG3KL8vToH3U4dHTsMtIskbyedtJTZW
PXHCiiGof/QcLnDI5DwqTvqrRUAu6zHYUBP5BhG5GsnznBvXCO5wJ1N/3tqyFjbYsJEUJa6LcKhr
w/c2Qn509rqM3agvv62h3RilKHrDkt/gV2dTQMPudy7BM9vBLcZemleHCM99/J8Lr8x9pPGxPXMQ
uX5V/khbrsPcKs0xzDoJVS42pCmN6idwyHPkrXUSlAUFKj45Pmca5N3bE20NLA3DLH4csScijai6
ltDyKDX5RsRE0bqvXAI68fqkoYaljVjcs+Ou7de+GNqdq6TqaTjNefH/iSE3BM6SWObTr/ufajaB
9xIeG/P815spWl0AVZi3yiWaI0bCebKxgjRRZhBhZE9xEjT8pVxH52ECEzwsJasyf8tzSaL/+ncr
AoHd6y0PCR8Rx0IbIlwAL5xDbAePhhkW6pXGikOTqO/sW7kB5TfAedDIH7pezh/aUZWg97mmjZwt
UusSIIgxhW1QwLKsHtKVQHazEwPd54C/DHqcQiNHHImhFn0fAULFbPK438gwU1xhdZnjuQriPOCF
Sn+r+4NVy28FH/KJish1R08LmTxPTkFj3u/Vi3BTENhyWMFb23WtR4JA5jlMkeA/F2HTCP39weOn
bI2BbC35iCCQnlYpbDRmKpnku7NpqvzmFFoUtnsxV67YbEB0Ic8DXjCtkc8HteCWYu8UTg7K4/9B
tG6KTQDoeh52tlaqXuMw/x283h2OnoMmakZLw+lUVY250M7oF8O0JFVp4v5c/fUFWVeIgwaehVUr
9cwI9IGfDfHPHqiXgM8YZF0KU1VTZ03Xf9oDBPJ1iiEWbhjO47UK6kH67UpZq5k/MHTNp/q4xmyL
yTXEuSzooi5b2Cjh0XSB/pUoKXdOpTNc2karxd8+NsS5d3OtZvypaxmkyw9aJyF5Q0NoP/Tq6lHW
M0A9iPCXtiR9Ab1RKYczOLPNpwqfFi9oJykpvP/nfyCPFJ0b5rsHAmiALy/1ek/+Snat7eQbS3NE
SL1IvgeT3pfG8oSVCUVHyPjaMQPTqLE0G1l9avDGrLJHmoeMa5EjXKUwS75mkGvmcuzejAece/1/
WKPaSNVvVRt72JFpsRP/+GNUYy9hzZmyscooxSYhcgpUasv/QG4jDhI3qtFRlL4VH9AEMQCY7Sak
+zSB034MnQc2Ekxzy2P9zwK6+0Kp6wZfSaB4+xzxu9kEwiaZpdS4ie9FNHLtX5D7fbhYMPGcRc7C
zB55+iM3Qt+6K5ypZj6eDLrWYUTT3w2wx4YpPx/fycaSMKOt1dv1H1aL1UQVjaCnfZB/YK+Z90BX
c3T+vOuyJMQOZSNF1IuFM5y4iB0WQA0Slgg5cNjSEKYqCQJZX9GZ4YZTrB9tAt/GPkIoMBNqN5J1
QcjAfjsHN8MwXKgnr0qJWnFL+xM1pf9Xtf7fsNOr3LMFn1kqZNuUnonaV/Mn02IqcL7+nVF3xIP6
908a91OXvIzFpC/FbRaqUS18ElvWLotD93oeNINl6L2ype0K0zfAoyJWh6x23RGOwmp3goHyqbb8
0R0I1YUpsm+FSFyVn0DKBwTRZIYrciDxxgg3Z/1qBz/20F7M36DI2SPOioZgYyJVXoTT0+hI5P0l
KOtSA7ckEw3NGQLrpWb6w06vzu3Jw+RRmusgdDmu23ZWB8xRwhKWo8KlnUb/8qcs/uhXvrE5b9Ez
jf49vz4EtPXk/BG0kX4NO0T/VDZW3HSaBE1eLqgeXo5xlTC3W06mGFiyDJobdoslrxNZEWsPxjQg
y2E4MLG/zR0Se6fk4WbpLedrjNqadruWCD7lmpiD39lwUg3oCP1uneDzE5xpyM1oEMhnYdEADMAe
H+uAs3NJg1c6eimDLEe86N3KTlSWnw29OMEfy3lUi7YOwL5l0bn/XaQ8ZKeP9XyCdeiEe2XzBYhq
q1YB84KbivJTRH/yj8ku3mAR6dd6LaBQlhWiJFlbNQ4h2AXX+g2uuqDTJyQTekTnGgDTZ+C7gAXq
yBtu2vUIDDEY83sJYaUA0hVcqzt1OWOAINo9FZdkBuWoEDaB2ZNVJUB59Q8fCmhoKem24mkYibwx
zMTj8yVJYIs+nIkS7/N5iIojta6GAnQiRMHEL4MdcbrW+uNwHzLe7Bh+5KekVH1WuPdtf3q47V7l
gBA6kTLEucI4PO40XHl8obeI2u/teUGTZCewBybm2bgKmCg3PVbPgMFAfLugChOPcLS0JouABz7Y
D0Hku6m2H693oE784/3OU3qOpUzWz9eESMJrdM8kPyUzjhc7sbdpamTmlhhfrt2PU6mtatWDPEB4
+bp4+dzyPnQSUo5t5SDqYQSRSzpoLt9lvaIAaHYAblhSfDmWIuAp9SQ4MSMp+OatSYCi/pINmFYS
jUvpcb8QRY7nU4nvgjH+OMG9HkzNJ4Gv151/DQNl57cpfIj4wrxrwPtOEcfTI7U7zBDU/ovkHCDY
XYL2zK90VCV5PnEFS+iZ/funt72ExNPvup03OWh2iVZ3a/ierz3KduEh1Quv6hwbCvRAQZz5BaOd
wGlvnQv4i5bww9CC+a13ssq5cZznrP332S7V0kX3g34r04zmITfL6NOFMudFGhe62XvIBkhSNpsK
ua9ElMsJqmLIXAkeYUNfyHbPfiPjLNILBvxaKTcZxaml4M88v/Nm754YFxj1u3Mz7JoH5iTK1yLB
zRyilqquUupE1L1QgtweqCpbdjf6FnwE8xfOPrP7sm4gtxvXs1gdK8eLhz7WjshoGSCstkNgtZ6/
BVQ8ItFFEP1PFkq0sgWThAEE7mqEb04Hczsg13umogeKELUd7O2c0smbMRx02npa2SbMCM8uJs/G
oxQnX9JPAVOFIFL2v0mUKpN3yYiPv6I/I6c6NfzjSbqM2BYx08mHgr+2CiLTm5+JdGUbzMQAkiU5
sqbBoYYGN6DWu0r4+ykHer8AgvNZzrzXLVuswg9Ky3Ktagmznx9VZu3+mSVW7G/fMJ0KxDdf03G5
DlEozjBIXh3q7Ra3mn1eFwthjnZddKO89hooLXNmohogJnXDR0jaUVwV0NnfmnQfmOo0AmtvOYMv
+bpEuM2XayDsERRAgWKBGPip+EEkhsZmmtlacJLH2u6Q+jEv1OogxP3dCu7W8CmccXKHQomSS9fr
Q8fumiLrJcLZgu0Q7gZHl4UtNTTmRwi5DtH33GekOyvc1mXZyHTwnEH7QCITk1Sq15P4D1YULJ9U
+VTLlpey2GjKUhZRX4qJKKrg/o2ixCm2U6bgQx1eByjEy/QV/ZQfrJ46VQZcSE2tb9mz0GiqN9PX
SBmynQKdBxub09UAqv1z5Rk57+7CNpvyVbRtL4m4/Si38+iejqul148quV8HRV5vu3nK6t6TUiNr
tG4A3rz2HmFaMXn1aYtM8dr01wjtxLm4VWdkx9EU74AR568jPUI7Diyjhr9C49BVdPG5+ptLCAyF
nZjur/pNypnBHH2SBAXQPugTdnH6CBvF2v6rbGV35EVqEgnffUjYSWQbgMEDE8NsMgLzPqglteRw
iYZRR/RxS6KPyFWNtJkah+jJ5PAjo59MSdgmXzi1WOQO+HwWk1ZCEbdQsFr4V85uBBUHq8FT+eh1
9eRWvGkHwyANPx1ov5S9VcCdTp2dJj4EoRbL5DNnCE1cqFkM6w44Bc1nbzaYLJYIqcVRefvCbEbB
RJVhKbJWKG1RYzQuuzL8xopHPBo31hCnZM3ekjklQDzLWSbL0ikYbBcF0uYXm2QN6J4UfJVuojbf
rfmeitGYoicquwRjtUQ5NgI+8KX9gp/Pnuvw6h8Qs1rZdtL4SvpcRmg16uHCocd+6b45NsVtqjhW
Gzi3o5o5nRGpzp/f3efB5VtkBuwfH9FQbjgN0vmyE7hXk30mDc0fwc1/y9pgaJA6/Ys7IiR6DttI
52HBkaOxZ5P1g5O0yfEcIK1CImm2TNKHn+heRhJ7xT5jU8wI7qJBkTsGy0PFU3WFkUo6SnAdyWxG
FQkS+1FkV5/KV84uvnj7TElj1oVuKSZ63XUlThc4AMstw3xS8F/3ncQZKbCBtEEk0RSt25cVPGKR
JMqoB0vT6nUb4O8m926fck8D02hH4UegNXazgdX5cN3Q3RsQ/QQxd1+QpZ7llieLORPbp71/jgUM
O9Mh2PP4Pe2J2GbQmxfxJUQjAh5qrNW1NusYJXnTrbrsrqm2yrFjmyjd14Hr7SmE7chOwy2b+udW
OMtogcRPoD55YjEGd4LQdkn8g4xALgGpEneSaoEBbmfBK4gbRnGYK/AotZtxJl0cF5Mbe9aRMWzp
EFHjhbjflRs/lDf2YECwrxGXV/D8CZNqWov0R3SKsXHDNFamHbAmdBWW6OnjWdp2oF0e7ilQ6NHj
Ae5wumxBPEQA2DTI2lQFewBbsMnST2IgBUdPANZNUidHOein/A1ZrcsRiDlFFrr63DrvhGuUE8z3
9y979Hjz9/xO9SBTRgnn2Fqzp2qYCV9v7+wIoJI07un4/hSsOchk0G+xcASclu+stFIrps7jK3Tj
8U/PYZ4bfnSDiXhAf1UUbtW4P2ip/4lnCDcK7qbDXnL/X93ISEsBG9kRLWJWG9NAa5vCFMa+K1wl
6lBdgoBrmH/CZyu3EJ7Qlud/HyyB3ZOByyXwyeDE6zpWqoMHSDG0Rv04K2AHXKHpP2gvYE6jH2md
O2O6N/Eziqqg2Bzn9A8/GpR0hEAQ7Z+27OrdIUnZwKXBy946DzPSvW1gP3RjsxJBtdm7HfSakys/
E+idI3PGBqdA6upWohZ+nYvYpVJJiPbrwjQBy7Hxl5c2Q6N2PipBCVAMgVfgv4ZoH9i6GMWXPbHM
ysMZaLsQeMyLe+6S+GHtTzLbpuSaAGBnq0lp3r0/i8wLjVIOdlO+u71wdJFZiVduhzB4IZp5uJm6
bWyzHY0rSl88Ne1l9Bc9CukJ+YKy+vbB1azrawt9A29LFRCqja6uznKgeF8eG2br05JULH2acddY
7PDiVYrd1xyKS0YbnYkwjvWQ/lUTul+xT2M5N3ixDU1nBOK1F5COwaxp14X5VDHfNrqtedpaxmyc
U+/5HvUztVcadcW6FYzNUdz4cey96pTuPM93BYfjaCGmTdbBoPqPExyEeqqjvIt+kwFBABByVx6M
ESe7x5tgCckXH0suss0pESAR1m0a0psVVD1sSvJD4RHPjh8CIX+B3uKdfJO8f5wkJsxR6HYvAAJp
Q99WNtnUP9XXQYPC2ZCxs+m/BumAXcv9NVWmV35fa3eey8wMrA/yn7FCgvQXvccaraWshVID4UDm
5XoybNQ6cVPQhsBXmFY1A++bpPJZCbiKle+k7hVLkKiv4j5bgWXxCuU73xyaXkZ5/6fDBddi6IsD
Iuc1rwlqSxspTWfS8Xq0Zcfk8/pDEQ7fFLJdEPP8h6g5Dvu8i3idT8bg6iqvY9A0ryqnNXfNnZL5
2sSV/X+L77Uk1vgUxKq65YuVaArwql13lN/nlG+XiW+zhK44HeTJfxyb7YtU4n/XE+P/VbCaJa6r
s8Rpjssx6bxqShv/XmsIKvvV6ge3hRy0QphXuQ0P1ve8F3gAWfzwRZhFP5rws4y0mHnIfqS5tw0a
ascEEqpU0icwzrQJTWcI4Y717qxUAQum2Az84t8vZU6JgFUhMf4CFdBeUDjMJZIEVexkP7RdaSiy
AHFyLTQvNGTBPrMLLLgH7i9wK4hCrbJgh0UqOt0unyLRPJX1us4ZC6Wsq/2nIgmJ47+h66JJka0c
S3cLZGsNomtNF0bSLoj/OOUUXAXW8NMnE5CdMByq2rRvhQ/dUvQKO/AnbhlwUymGkspMMjM7+iD1
Kj/zgZvo3O8viHJO91e/J9ByRqJG7RBukUOH2wAY8Lg0c2lfg0qnTJKe7PcbWTu+7G9MuhxXym46
HrHvm9zhX+0KpXIuIMe3g7X/BcBAA/g2W5U182ryocD94+LofnqyVo1QaiLSwK7VGfCMMIIHXpBR
YXW0TUuMnoYrjLN9GNqLxDdhDBYIzqheQ2gOQa9BU7vGcup4TuCL9e/QaJWOQUTr4JBxXUjNBaMn
qaifAXzp4dFoZDPAA8zTKngbcz28uJmzcXzakotQP+qVZxfKa6YfCBBgOjbDta3+W6ZEkUZVUKmc
GX4aRL+aYXOnlyoeL7e18aNMpB8dDUiAf7zg/moIrWHYMJoGCG7ZPgl9ig1LJ1ZVFnG33k1y4LN8
SghXvvAfMYjG9JEF74ebZh9X0Ka95b50hm1k6+BlPw1psGCMFYe1eps/981NwCF+NzygKIkLnx9X
NUPl3n8f7NnpJjVVrio8Q7wZ97LBNG5kwtK7xx/+p47ZKXfBVwH++NojwRMYGXY/YULoSmO8hfVy
zJNceNzHq3AaLlhpZyTFMCRSJF/OLEQRC0niBFNf4lra6N0CFqzYfx+N5L7SRgurjQlGOLZ91hZi
IV0SGkJ7XERV9IUMcJ8TZ96YHcyyNpE1RhDwxImjdHtOfobjhxt+v89jRVKoEZdFz0ChvWqf5A8A
6UNYXupwnYsvq++k6+YobHAfAvRZkQbO2OLksbBk0qjgnXu4YlGfhEXvfyq1bK8opuP7OaHWwDde
fecLSfFN1TWs3ZlodCiE/6fCa+lzlaUUOupi6DHGMIlc/blXeUOkBoQxtaAgznUOklkDy0o8MjsM
oi+bfp+Sw8sQdTC/oiV5LXMd+SmmQEQ1rAUDTbpZPsKoTJLnpj1FWutgdeH6dGWeK/xXvFciasxw
5RFpj7d77GG1E8G8r3ptD9z9ikIIEjzXNi/1qGyFQHe5jyWGgwumJKlvXqNV/BOgsPf7ecAX8X2q
meSpe27lH+RDZqZ82nLA13pMl7/7xvzv3jFNCkLKY7YHMXRWKZk6wQDm0QuNWBhobUlOFqrW23+C
sb3t7etwyEl3t5pTHwKEuPeM+9sCiR6BVQ2S1rVAK/WrBhteWW1hWDEqbYGUgQzQob4tCrNCiPzc
V5dEvgcqcBSOii1Gf2g48wKsiWtyiEZtQjPcpgfKp7UYc91QiVyw1//EshNdxRp9HtXyxHaKKz09
rbKSEB5FKPsMjx01jnWlN5+RTqyM+4glMO2LJIF+vH/Z/cyKbmyMVk/4iEdHFONfYEfhtCmCgm7m
BxmQLo+B4sCjSNmxxQbMCBtpy9L1lOH0y0sUFozwUryIL5/rdbACqEgUM10X5UmXVuFSkNMp7Xwi
La04g+L1/TI/cS5D6F0xP9Eq8IUKaNaegizyD65vEDlSYvp6j1ij1kVOwuw485DMx02jgs7Bf2NY
OOa/70mLJI4pXlpOlmjSE36OVR5izuLXAwqnBQfY/Sh9Dn5eGw2rvywjJyJLv4MJOBS21krlQpVn
gmMC776F1WT5KrdAa0FRs2QAs9TSKmxnc1+DD3i4ckNcYbAl+DFiJS5/dEmobiyDdhLqIV3McfV4
fcg7U/Hzl683+7NAFbLhfx+8dGU8DVcsgaAZCefbTPrP4TYLYX0Zo/5YSwKf4+gsvsSbYTTLrCeV
5M2Ar6w1PybgMegdIJVuHZ8ulPXN0FNSejOEWsPf1SThpFP4OTvfo78srCoBNvj+SXZ+/a7i4txm
5wUEAMuTPU2MKZrv+zm1u7xXgSTEXGp/QmeOZK3mPtc3GKnHy4LC5ZA4UZo/f/C8KjwwmgDwEtyH
V9sPLLMB3rEF5N8uLFBxWd+GRgBKJyo42fr1D1Qxu68COmd2yVFBZL7T1S3rgun4MelHv9Hsyn5N
MR1oxncwSz2v7vyryKFBTesDJJHK/CtgxMbfs84XMtwqSg0MNrVD/6NmKQf6gEFQXW7/KourVi2h
gbhCwwJ9FvPkZ5lCsNiU/1FS8XBZ66RyIGrwXKs2IJpGT67HlOfRGJEML6kgmkk5mx2+0uf1EuBB
refN5m6+3A3LtXXcE7Hb0GqV9SXwyKW+l8i7+gLmYUxTRPEZiXmHeWj4dAng3OpP1mVLeTXskOfm
bYaK436SmZ6Xej/dqdTu0t915O5MYbM15+EisA2yF+5nC+HbQfY89b4+F0lpxBWQfSFORQKYxH0J
HfdeMUqPnthcJSxnIjIejnn9gVX++2U3hOAALKOCz92PJVwP5WAIRrq6JB9A/eT5eoyja/TOYifp
EEOBf07fQt5VEQrSsGizxeQOR4zIkrC2x68Yc5hvZXHQiv47xS/qNDIUMsGB/irJzDPyY+dg8Pjk
kQR/RgmBxse5eTcqJGPCUbWP+NUbnN454xhQpuk0UN/8SGjCaOx0Ww4Ug1BDiQ1mSKoPTSuCQLr2
f19goKTfZtJSxPxvhLjGJS+FHFZ4/6kpS7Vr+LdVNESI5tITHsGFwCpeR+rZhH8a0KhySfmId4/9
PFUdhGjhTW3FXepLvpnPFz7c2000HOBekA1rZbX0V070QfhrRFFhiGWDjN08TaVnulWM6hUkxdBI
+XVMnEbsdIq7G5scC/rKjhnDX756KgMDoK+3CYyhnHVaDqlHL7g7hrMChnQLLqctWRC6n6i7Aq4v
xEWMt15BeTUKruggY/OMryUE3XMyZOUDvMTt4Qo+12aa1Zx1fJzuCI6vc8ztdTYgdmhH3fM3aMz/
93hnTbKvdbwfy+KtlvK/rLF2WACaQwUbhv+GPrqq5/XZ8sNFOYxXyN4jmKLr9Eo24IXKfbK+hMRx
3ZmPttBxN0gL37pstoEqM1m/aL5EKiz79J7jGsjLuZP4QhrQCMB9lQ1xzuEBrRXVm+iezJlD1G8T
cLlFgoKDNp+ULyCLCQSUof6YalK/OzPpuoRw6+CB11P42X48vCbsWY23zQPGWXwiF6D0oEtacDW/
IIu5P6FZ03zoGcrL8LMHJNlugCv/3xHXiA+fMqC8qGaXgq4VCSBz67GQzztQsFXLAkxq7Lo/5NjM
H6pjY8baLndLHHEPM4EF5gTguNcniJwRXnx0q31y4pRcF4YzT9LV0+RzMSQcpQZouneajdQtRq5p
Q2mhmNUPnm4d8IstNPa9FTPipgDHJzUrwFkxdO2MSRQHxdogtoLRh116TXMa4OVlw/a3K6dyuo9r
m6V1ilE3DRqXFNn4FVl5cZdfQbYzkmTUgoT3ZJGzbnfdVQiteO9x6BCECe485ddeDyR8eUOGa8Rn
mrcNBx8RU9ChMCMU1oix3J2I0ENYAK55FRN7vDQnWJceU6gjAyYhkZ1XmQX8n/c4gAgaUA6FFar5
kyAmesfjZzqL7++6tmBizbYTbrg93zkr2HGEuC61hdZK1h+YOPbnK2wd1QtM1NYSm/nqzaK9OF6o
QZuqF1e2dfbKLhu8bGGjLDLvrwiooyoED0xURb7UrZbFLwkvgmH/nLeWpzxgpIgzvlhc23h/Z3jr
9atJCqqReDIkGKrG9fxKLAgJrA/TKgkj8ljfc9YVUONcWBFWo+iuLs/+R5lpHqrDk/qa4aUqaAXT
E5W3MXZ91xmJH4YuJSc1ohcaEGDAF4L48MBUGwWncOt1CeopL6jqWbZTTp/aZP9W47aIBBRyC1OA
jL0Vrkwn60Dkt5PMQU+0JS/LiVrqtfhoTdmN+Et2fOkH8KC6DcT2ierZIloI37mBvRYppB/TXXPw
IFF1IVIZx0eZn/WTOYTJtslsjQ6M7C+lk8rrO5pMwYZjP6gvqXDPMa6rnnxacYn7IEn9oDQsVUjE
n8AGt1pJEZbTLa3jkWr6/0VEg6cBuM5rmErlA+lNmyHYt3zzqBD040L+AgflQyp4lazWGjIbyMy3
WMHxZ4sW63yTjFY8DmcPm9CjIUfSQje4BcgPYLrk+JfQjaCbBqmCw4F37yWnjfDeMbkoIEvxdaxv
55iW7LlThXgQoMtRGqd6dVPSGehicFgDjsstGJLHjon2YO0UNKJaVeGwEo/DiH10+Gr93xGAyc2k
9e102BhItaVoLh3WOV+06SeyNjw6/favYis/akJjYNwfnUHxnWI/xo8DCHkSedPEW5LxJaAK2D5T
3Po7YkhPquA7wylsNz4reY5vZIBfl1pJ9plsAG8adZoelr4YtEZLsNp7Hf6x9fXhGJZN0OxGda3U
d+tYX2SohnRf+FpNcRk9i57nZeFGyinNGR9jJDL4UL3tsaw1f4ILIskbtx2Vm615oNJOY0BHZLAS
OlrAXM4Q7UiRps/XsguJo9NyYIGbgn/7sWdKp1mk/dhb1/riOMChvEAKl/Ocp2ya/uQWsqYtGPzq
N86E7TQU3W3GzdePgqDLf8YJVCEUtAtYNp6scJKBmiGMnHSe/9TW/1NiL0VeILd2OweV7oXnVUYc
z2vyRVKXykzhIzMMFFVVpNmsbV43CsFXA+BpkRwQDFct9xq7jS7V/2Q961oQYyzXw7hKvCmUaD6z
TGyhGNA29eiAnAQIKBSTpj9r+VobFOHENW2HPbMJV03WRaOT8QcoBR0E+Ks7fQH7thEFI6J8mp8p
PnFH+SNMv6/PDW4P/ZGap4xIYFt72sifc8/nsZAbvBjOkt4+0vwXR4G6PrpV4HywFAHWtfle5LIQ
HUmI9QViS8yo05qx8CMh83bVMhzn90XHGYTmIf3bz0hV547aylqSgDx33khjvXlNTpBDanvhdCVM
QlxJcS1TDBSyFnAWOemhecmK2kKGsfKC2qGo5W44Fx6EzBoPQ4NnuaC3M54FMx6R+mh3mQaayP1o
8HMa4E5rrueS2iUm+x8+8lMWW5+0/Nei8mEb56Csbpm4xti//VMlWIxmWv/78L8QDaaSY1PCOX+r
bF20lJleYTJ4XnwQ5K/qsQUBcfUt3xcKIQnUJ6102aj1fLbz59hlvoJ97Lv2+nmS4TGZbikYoBc0
Ol1d+GU0HoKLQKKNupUMY2YbqfS4NQ+hD/Wns75FCPDvg+KNcMjowADc/Zwp6lTcUjNX74OBlbGI
9q8BxxSH1JJFzTruaNZuiLLtEbakstEuhB6eGiWRgvmWEssIqtlNF6wys8lSRTrdYBKlFqXtpZ5W
jQ9Ojwb2uVWZkBEyUDiRhKCB/Gb7qqcWbwQhgqPYOvK4bfzP0cSyo9oazB8o3rf9lrc6bEqPCfwZ
pB3Hh65Hycvm3T9nKRMBfhPzPXKh5cpvLOiuMV6o7IlEgGeg+8pJnw42e5t3IRx4yO08LRAIJu//
7jXTCAVXpsWnkYCB0VR/EFbbXbLDziRn0Lfh5KFfis913bR8RsWBrwetyrbS/cVgDnRkpSPfTebP
NAEg1LqhHYDO9rLhYS1pZw9oZCq1NJvHbfqcMrni+ESW0jLWlQPQr2kzb+8CwTLTkpQc0S56iu+H
VkIrKwAtb4f0PC+QlQCR3QrZhYxi2Y3UD2cM4zXw7I6f+mLo8/whpA/8QRiohUf+Fw3sSz90NZtS
C8dgdwIGf+O67cngI8dV3yvYZZ9c5ScbJqz5rXJIpgsD4x5fsxpy0fuiMxu1T2u1cvVMSdmRYIZM
mj7RX+7vvbIHjJjvbOzo1PH4QpveF4vssqTH/HkL4v6V8wRhzDxPzCiL08+2jdaSDspT2RO439JZ
zuFm+aoCvFijjav7MLOC0fzaGWQgoG93im9Qf2bbkKS1XP0qKdFitSscLL/FB4qL/LZsi+9CZ2bY
LXUVxcVR5oFRIZtjjmQdrdeEz0c1S1Q19n59oTJHr+L9b6tTrG3N1jvIVmppdXwq6kgFZ1+GKCGQ
SmCMslrEkR+0VEBhwvQ1TZHrQdi3mHoozzRIbZXsWrx6niU/fklT7xFyHYxD2/Z/+aimlbi5okaN
PHTAr7NvRRD3LgQ8mdAx0HeGCoJ9iaQAeM2cnp7xdhaM38w5VbpEqHwUCjkgHNBYntnl9K0nSbs6
YRYAdDKTteKKrOGYiUpnZO15kB2Wnc1dj15vXpKW+jnaKN2C1we2aanzWlX46h/aR/1CK8gyOzPB
56/sHIm+gbzs4udQvoBT5fPUV+pOO9S2wn8QaeOm99BfkkXjrVNfJejH3M1Z8mEhgYaMuR9T2jyy
MJ5wbHRTVthQoGLu73myA/n8rKgpPdC8LVkdYluwhEi5Y/sq7KNwlaGq3NbO2SwwFymKGY8yNn02
W+h6fLaUh7tAoA488rBDnx7qSO4vnMXSg6QuB4WRANqnr2bPLtwFJNElwhhaD3qplZ0yY/Mw40WM
EB1eLPC9n3wr74SJuY1MFlbqGk7l0pW1PMn4nxQjW2gx/uLtSQU6re4nAlO+cMKcpmvxAAiVF9Oo
K1Tk21b9thzxxrt1GzXPjJnAXOj9HyJSM2BuNedkatNkUlTSstMIoEnJ1L27KCJu8Ww9o3Y6XB4E
buaDOTcfXc17AY5JboKH+79hotPw9pbDBcjhS+M80U4FQPQtt1pcz2bPVWuexWpa07xmZcCUW+d0
IAVwapiVKEAK4oeVvH+T1rpc4tP8Mnp8sEIF6NdxVm6zzeYERoAWXUgKuAhAW20jivY7lY4luX0m
ygV2lWaI+Jh9L28J9CkDSfdF+d2eJ9EU+KalbK5k6e1FtZoKiQxWlaPeNg2fXpxqv15wgMXniWjp
DwyZbHjtgbV5UxW+mTC2khlx0KgxFGNKen5V3ZDtk8NMcy58nzCKo782NS6gLOMun2C/efReyahB
Liu7hqydBDlmaVB62lnXLG06mdBIGVXRNoFEEjnIsY7W9eCSpuAWhO7Ca6sUU6ld7FQb45pnYkDi
Szmp09SPRg0x+tzc3c7iTzkiJ1AsowkgGTiPR7g36iuocJDPaRgoAIDBsQ8+XAVnchSO0YlD4+Pi
l2Nqfk1UhWiNmOVt2Qoulxnucca5KPMvYDrZckZEjXLre+B9gh6SIIU8wFCezQ+fjZrC2Hqph4u+
y/DiUpOYkPwfXpL9KbzxAYMJulc9BNavquiJDt3MkT1CLCNK+kTkG2a8H2uzqsy8wZgkJlumiL2H
emWjgloXbl6DBweu+YUlhPUvvmxo5Zhz2EK8XampZQiGiPWtmqs172uqBgirtjCWm87fkO6AwleY
yu4lN7UwT/za9z/hjDvv6LZLWXhA8qjREPzFcug6ytgXvlDNA6TUA77lSY88r//fMMW33GPAvK59
Vd7jNuEFT5nl9V+5qjFPhWyh3o194JX+74X+MYUyY5Cr+yZZBWqhEAe5Lpv1wR9+Mv6kp8gOHMgU
SecKKs6sT90GN8kfityQulCVkM88cLNTTXDmthhXhuOcwbL6g00n+gnaSwx1szjewSnYPonJ6AUQ
sZOh2rN2nM67NwJGHpG5DIb1wkXHMdqSqDjyqgFSyWR8JVNsR2VYn7M9y6+cEx4k/pd71R9eqD5B
3zwo/tDUu2uQFBgbuESmajqubr6HbxdAgJRPf6cVuphQNQdK8DC3h8PJWZSgF8xU67xYB6HaPV+y
JnEKQ+ZKi52YK4sz1aB9AhntAA2p2zm5S6Mh6MA3c1U6VZkCcpU6V/GH/fgWGZryR0iT22nB5CNu
drypoyz700gkNn2fTAanjDodIyvv3YBYq6GmN6agxcg6u+ksjZ/5MCU57ZVIAJMu25iA7o6pYf5L
ExtvUaYpBRjdVdpwmWQUvQreSOthDA6itN2Pv46X8e2Afl7N8BbVlmbJOMatY/l7QfeHYjFTYQfP
S8+Scj9H91kl7bmV7d77o0SwVaQYUGJkX0uqFSAAbiSiimSizdIn8h5Ec7v6n6fxhWVsO8eLsWQ1
5xpA+7KJjGXmJfjIZoDJSqNjQZPXJStBW52tmiUwNcjuUalYnrQQIqqC+HC26st7qSCfFfrzwtZ+
5GIjVsJxrfJQQihz7dTsCdBZOpapMbBFDQ4CE9iayWcmDXv9kEly2dWbemMVnnR0rE76zqmlloPM
39gUBFoufv2n/xFY7zK8YYg34rviboKMDvBF8Z5yIyC56DUZprO+rJrQEerbIrLCh4VRKf+pnrt+
14coC4QyXPgZLUA5ZNcmWqYv5+7c7nZE4h/oD38kyvtnmPQz2uj//QGee3y+zlMncu2vgpGiUB5w
Fv5DcPFxm1X2B9ViZY11ULKAFyutdDSjqKuQbzmT9vLClFn7uTxHIF00n7oeiSx667MK7dXq4DHG
9NBFqVVBrLJ390agt8tamJNRuJeGkVe2gHfH1mHyVwlRPBtg08EIbfPvyoZ5jLUCBFkI6Fdx5p39
Vup4py+RKlmNl+8zledo7FqTpQfz7B9m6N/wivfLX69M5fZpSLUyCI5KNDGfsTb8UAknc3ZI0YR9
dU0zG7ZX1uUSvmQLP5mqeojamxoTa/LCVHF6LdeKwMnNT8HwcPwauYJifqslfLZeyJtxAPF+NhCz
QwwGiqUO1V23vPkB5NAz4vqjExkucYbFs7TCAbHsVwv4bsBgjsfDGVd7FTvEuZ32apV1cz8AHTrS
YTFwpVuxiDOw47YvMpuRJudEtupJTnGvViVzvPwZ7xJrW+F9+Ea6KLWZEo8UUGqL+b8XoIKTgO/R
USbNRnLaUFa97dDBBxwPCG/lP1iIlSHUznSXotdI3RoImdbV8B7u3Kg6/C0WOScdyTCxj7P7iTb6
oQJKcfYMsacZJu6pAdbvVUO5BaWTlS1bpTVXZsbzX4RZ0EZTBwBQFcYNLL9vduL+gZyXailGUUJF
SNE0M2E/aJmhP2ZFQacyatB2fbL3GGBcA6nmg4EwQFubxHNhEQRyKyboKCfKB+0BmiPeP5QJma/G
uXSm1M4g+VYDWvXAkgpYA+Nhc82QjWFBfHnAgRs8hPtsct0XTh6E7slP0q6wdaAbGVWa/9UT5UWy
sjCRFmI49MitRXacn2RKAvxsnQRT9a09Ctv3u89XG13sqVVleHPRij8E23sVuYk0ErY+7fidQaTP
CMd4mZvGqGm5rOuoUOPZvo+PhBoqzEwpPU/w3Taj8d8d553qK/9WO3mP9Zw0cnhYEZDs/IQ7gMS4
pfgS+NX3KhxlhrAhnJu0zlmVaHojISXa3ts4NcSi/rT7xAevzBG20+MoynU8jpJo66r8W8cWtkgK
Eh2PexWxRA4bhLDupsTLVFbc+twIH1A7PU8fzaw+pQcZZzxGEioLGWjISS+XXR8+d5ELz2c8LKXc
7YCtJgPxxyj3soohJvimcV1ndvk1p9Q+LDJlIP0aCjNOfR+0KixSnwMf6sMj2ngkmDyDRp5dyY2X
LL0FRyiWoUZ2hmkUAMw1+IR5Uf87XfZaonlvClmfEFZampUguhGo6BZfaW42LUdpB6lqhzhrgSdZ
uVg03daILj0gBMQcSMyKu83IqEp/KBNiCpZJt/gOt3y+EqrsX/GHdARGjEjGQvnaaCrxlkA1eo5v
BGOy2OowTSUwdM0CTZloQ8t4BqMf7BTif/5g+sAZIBfiERPvzzM1BVCqSlT2J4DcDLlVtote3+uc
2uMbrwgq9sQiTXJahkv9qIwL0d81zpwfT6v50Cn0BVN7AagkkEEp26+I0jlyQq2mz1U2uCvCrxvY
HlAVol7z1IbxzOkDFQQMqNF47CwGPtkl23Po72lMbgCYHz4F+/HHQdBZkQCN8SM9YYod7pvpsRGW
h2TlLHPRkEanJVWzz89H0bLjyfI0jBmWJuciQQJBMEWzSQJged8U2bvNnVYY3oNtKNg/k9KweCSG
ezF+qCrmiM2NmsTJ9d97qMjS2XhlKc8BRJDR40ukIJrTvVQBR6N1hO2qxbEm0pViGW6GfNAcxMgD
Js9rtJs7vRAvkUfb8Se9VBWC4AW1WyA8LUz0ihb7iE/Yaw/hayBIfjQ3lPQfXIV5Sg7z/00QOins
rN2hOkUk2KLnKpJCSglqxsPaZwiX+OYFGB4BdkL1KI0Acpq65N48dwmgOYdjD8SIog9nxrT5mWEX
APR3J2XhUi0MvQphDtkRkPb0PMqCbsn3bbRWyKGNXNUa0UONNpucUYCT5HVwIr5Ds9Th+g4FY/Vx
b47sBSjgIshovAdEWiQKNXmsL+qbC2iph6uEw5iH02xlave71GnFh0fnl8TreIOGINta/cE1a42k
dAhFYd92euS60msGscL4rVT4QwhKw3f5MjgL62loYLH239rEIjBmbY79a2/LT+MMcEmfF2Ovgvf9
QHNvIdIx0PEw/1W1h96Oqf7R8kmETfM1mi+pgblahFEJIUVDGF6nqiV4b6XztQ+OXbQYFN/d1JvP
urAhIIJABPN5eckY1GE4hnF5VR06UDFB+a0UQbwtw52a31HOAKAywR8a986397gCh+PW6oqxwbHL
IArBZxldHqT4LC9WHPpXqGFaoFx3ZWw2gRX2UaHISryOLL85GjLOreVZywXg+foYXjt5SBsZSPaP
QWOS9Ubgv2epCFInsaAs2FqohkpVU0zlKiIiJxD9fwRSIldMAFa6YYb7ScSTCSR2H1IKWhtoworu
zRiKl2K8DBaZh8Y7jemFutOz88i2AzqTCux4mIYBgfSZyRhMd0ww/HwInI00KZYXfaXfbNYyH0dX
RgNHT2xjg/vugkme4SQcFgXVVZIcxsmgweIN6MPnjZpCsriPiRNvxZh2cgSaoPQCSaz/TVIGl2oW
+Dk4qP7FddZZ1bF3u5cUEMF5JtehmnWssvMr7llL3RpJFsYtjEKONgA246zo59eXPpEmgHncwviy
uphTISiBEO/aA5S2E7bMGsvh1STeIpsGgf/AsFtr7/PoskGQ8+85yu0xkKnTXsQAl6sv9jCByCQ0
VwE4hYJhZzqFu1LN5+sQp5X9gY27yhRDcTgMWldShrnBH3rao+wnSNAkkyvX/wqT4cFB8PBA6Cr4
HIwUMBdXYIH4gkJbHVzPck1FsTwGQ98lYpUUSRjsPnO4EslP8gBmbc/FLWJi1huFZTU2numTcgkM
cFwGqyU0hUEmlN2eL8VdrDqNEpoMcJV94YqKrO/SquOf1HdQOKwUwVndbdfB0JvOfeRo5KPuQ1wA
oERhiAsW0h8PnvVWU1Btph+1HKvROjr7M8E7LV8dKap/r56NgQJI+ZHusIXasavHvEGqKOE6T+dI
xCGmOa4BtRjSqeOyjkyZopPHWbq9Gjo+XIS93Tb5tE3EFdvVrce0tqK1yPabBpjZzFpB94wiM06n
fQXYYW3m8UCQSWdQyop6kwLXLEfLjVqj++D5/E79iNbk37jsUyPht2vF/H9w290MUP91W3GLjGu1
EPXKk/mbv/g1lOQ5HYoAN9CcJhH8BeHVnP5UaE6aPOBU7Ks5xAkbC0VDTvnDZI2kCeu3oxaz8pGm
q98oR49lhwBvVgS8Km8z7tDzfvWA1P0pJq3raxljNLpjRWczowG2UII07HhkJXLc3acj8Jcmwa5k
ixiYiuxuc5BIsWYNEAUwyUy3eKvD7ommtxnm8lsCYqdnng8QcUED5ruawbYGTIwNMCjo1bpLtTlD
z2nYZ7pjIwqSudDYmg89cv3PZ9AHePmP/MYj2P5d6xgD6/SmAZ+eRJOTMLXa+avECC7m+JgZFJbl
3CTQiJ/h7rzaA4J0k8Kdr6WsPvWWz/6e6xoFnjGKQma2cgGUYNEfbjw4FrSStnanvxm0yk0uluwm
o7oC09+8MUjUQmq5HqCJP9XZ8L4+TMaZ+NPQydJcDYat7uhkFjJPuV5ykkMiFO5ilLsyIWpT6DQG
y0UibB6pRmUcYlF+iz1/NZxD87xG2YvCCCPopAeNOfGP3HrzXh7kYViXpt5meKMlQvHW1rUQxoyM
G1iiM+FKt+U5kt6gcr1B5FR2zk21Cy5sG8KK0QKZFW3qu7ZluYqLrPwc8g7MyCr8i7wrl8CeZAwb
5za1KqGjpdU7j0+5NGggc1K0ovrSw7N/DzQEe2jZY0NrshDx2gL8wb7mcU49Nd3lK2rQErxEQpE+
JyrIJjfkSaRjmtjpw6FOexqKuekUxKQrGJ2wyPK+akubiOhZOPxqAw1wCEnvn4Qqx8u7LLZwKxZS
pLUxfZ8al15D8Syou7bbOZmBDnrWHQw9u7GUF5bK2HVtFmuJrkFuR4Ms2lGruyIiQcqWqnwSEgx1
rno3vUVI8V2DGK8wpwVjepanM0Tj75yShzCMr8DA4qv4xncYojSD2/oNkSLcVL57pBIJmN1syozM
9zn8ciA7BQHmPK7kDv3aBObryVY70HbBs9psU9Z4fR+l209lZjCwPq/4qUXsYFPmtif4NKGXO4qb
VDD0yV0geB9MWAg19s3uVHOF5ahrzsFci0g2+KuoLGt8m2/TRHNCthKGc+fqhugQY0Gduvp0bQBz
zyFdATUrUWf/WBy9HtdOSQmtvXSCvUvbC3N0tYoi8XQeUuPhVPXrZyvbZ+VhbmTt40f4ECuYP2Dn
YjjyyGplR8ALrm9+tEWt49Mi2x3ZkGaGVwGkSuA9ZqktmolA9YNzxKCrwubKh46lww86LaDhcAcT
GB98Kx0NpB+n2c40WFur87s7QEAuc1M0ma5H3NlfhZlCDEpr2SfL1itTbZmdNczEk6BCOE5gyha+
NKo/mBItQjL0YHc8sbEZvHxiKq86R360zQIHami358fgLVHxqvVPyAUBlT1w6S7gNiDWw8MoHBFe
XrPkYgSTrlIiEo9WxxLHdjEGZCRk0MdrVZyo0i8BAJRo/33jeQVF3lJNDtMwgaQT6+x/rXjrxXS9
McVG90qDqPThN1dDxSr90w/AO8CsHuPBlLjW5CvUeT7gQSEgp3F/3bdeHkhdwM/8H0MospsUJv0t
uYzHnsn3O9WUH+knO2oOAy5J2Z647Hxz3s8CT/oyfE33UZAmWZUySWs5H+NWIn0AmsXUflX73XbI
nyy0HbLFxoqJxnlcQMwoiOlq37oLCZEVyXTM8InUhKTp/PBYcD+Sbx7pVDbM1BFPM3gxqQFbpaXa
dKB7flLY/+TbsVAyOWFrr0ZwIbKG6BvchN+GBkLbWawwh+EHsXAzztvxXfHFSDw0CyQZw5eBsOxH
jCJwqqrp69NbcUwzYfu70xXogjJg/sZOXNM2XcH1R1sAvDqJCq85DfUnqyy/npjzzrLeuQpr+H8q
TRe31xrq42r3DSZetn3ySftRX9Dv054MeUNc9FO3TLo/Ttr6Rz2AfrMNpYGxsE2U7WauMm6QVBFY
HzUFkMBV1ljN1cUVCD4S5V39w7BfL4yRkFWDTgL6G6ro/eVNKyjJzyKZ9g5ivad9f9eMhDQ3/amg
DNrKMlRlfXeN3BhSeIwGexjREGIUc86mjjvFd64b8BJttn3TECEqlqgGNrvXLztqy8xlujkM8h5N
l+6n31awh02O5S2RUjQbFuKAvbL6V4OHDoGbgjbGnuj1aLmMei9pdc31nuoBSojB0pFVNowf7GCC
mqTX3wf4Nt7SvlMLsztamasTuXSk5y+n9lfNHSUU8sCXVKRy4TQZpld58prm4WnKc3mUmY8T8HO1
K8MPDYar+T0FnSBkrOTqh7ZTxa+VmAfom40jAlM4vDR369S6eIN5rfyC6dq6vv/VcQABi+45lMy3
L3ccfSOjszOMson3smX3aw9gk5vA9iBN9INcWK6sbBVHPmTZy/YO2pZC53wy9D7OrnW4bWEDvuFB
pE57bGYstbkvixBGoA8iThuOPZzwjwYQXIi/QsnxIKZOpHJ/KXO40umz4N7rs6oeEU0SLvqgQOK4
PYI8BtE19wi1tKZE8ZVQgdOClNpIgJwEMRtfy8tBs0NF+p+KtET1dlnQW4/F//3lrxWnWdWy8aEf
xu/ECHWVUoHLC1F68Ru/2aGXHn9ZbL10uLxHtXT9a81wL4nlWKZUjLWh8J2hzw3r+dQruHMle//m
3lX6eW0RyJPWnF0YSAY/wTcvKhMjP6n9IqQRUIJDvPJsyQ0mdRnTObTL7Sa2CLgE1xPI0Ig5YrLc
JWZ6FUqJXBtp26c647l4ZfbRbBwHTMdOi+5yBRiYccLmH7lcHQlzd63jvpBfArdWA0Vj/1vcOumW
5n1qFoYNO5h307Vq01SlH1XwpzwmqxD9Ocex9H6VzDxddMDAtGoCnLjmdHDBtMNEr/YTsa8wAkz2
YPMVfomNmjrwczIgIid0ocIfKi3ErnY7O1DIOECdcXEj/A7w76nlbEBme42YOq9IdzV+NrzpyibJ
vx7flRfec7zF2nawi/Q1rHqf2a7l2BEwmXdLT2mXuZNSOflW313hb1yKq0zntdpO2c2xsbsaGt1d
rpy9hu3ZOsyIcOXQ++tXCbyrROJFGLS1R4RdjtoQ9gTfnouWPXpEqXQjqdQFunoAz6vfC18OeNnz
EVmhCodvhvKXtwh1oeszzGPJrgDUD15gE5NhmlLvSbc3y7v1tFuTcfLCfWSwduDbPPzHNt3zrWQA
XvXI4WNzGStcn0H0zKEtdrIVElPJH13ntgpZL1UJVHXpay9weF6cd88c2gBDutnHcrJ4O8CbU1/k
4zEPJpqjULqWjMx+vUS+Sj4/pRENt0PyBXtcJszhFFrTZmndAQvLbrlj4BOfqV0RMY1V+NyOOzc/
iBmVTz/2UAcyc2FMz6K39Xeod95A4lXytwzVJ0g7UzirMTw5FZ1VDZu/qTvFQTfJ3Z6ilQnddnFn
khs6Do29lib1BOW7oYk0dA93DmN5JgkXQ5ZLom/la3fAr0ubZrHHGqWHriw+PNWzw++k3dj2c/FJ
RjZ2cpcPSkDGqRFqoTmHGvzJNr2mEHEXDh9K5VutrSOwS7rgfKWGGvA2c5xbs8rSVKRy4YP20jDU
j8JJ+Fj5yBQ03qKJeFucwQ5JHfbfYazGQ6XQf6bBT2+y3soNjrjrKxqeozx1DhGrkrhng/SSkTGW
oKWDwffou47rgy5WKKj8/NFCLwUTc+MhiwdhnvlUwbF6sP2tr7IqratDKsftuUPkaC76IT8lGv8I
ysTLvKRglg1fiRKpc07nbDbZkjE7KrcBcSrlTo61b1PnQIV5y9tXeMexlqTnBUkavC2J0yUc2uUb
NMWgG7Gt7KZo7w2FBrij5oktKWFaCGJS2ULFhWDMb9TTi0Ykd7cTuZdQl9gx6fq78Wg/gxte64MA
1Jqk/mgFbg1VoObj1EC/I2132kXpQEvJk0wcXmt/VHNjcgU4Q09SyR5WKqSD6j5/DZKKQgEUPVXs
VdmvfiG+0pkerIuf2VLNQAmpxIoA5N37qZo/M1T6TMSKIG3sIf7D6CQtzBx6SER5DTG4K1T7gRs3
3m5Tft0bk+ryaQExA25PzIrfxN62OPCyiNVfOK/zvDHhqujAWwkSF2Hb/ta2Ar8pkdp2/qLlQi/h
lrQM8uyC6f79gCZgVnuVUxhY1KMRl+1PA/vVRtqNcnMhlDy9HYiHkN86UTer1uD7lA+pSd4382/+
qPfALWqYBVpl8II3+I387qf/Raewy75FVk1Lm/DEI+Dt//aTCjjWylc2nkdGZqPGoowSSk0U7MH5
0zkUZLsFWPGJ+cuaLctmJFG2gX78OUIxpPmOO/YSOHABdRDTpGO0nDTcXsp4/xSXJ87VfVwizZ8a
L1k26pWSMqbkrPW28rCdmNmF3E1vN0fj6qQzjB2HD/QBqZVAt0gYEAb3w5aIMi2o3nL/wKQqRhFr
yxmyd7DGPawVAiJoSdbwq1tU+QyNKNMeg4SHc1USgftH39CNj1p83o6AAQK8kvqcZQ7lLDeS4fEm
Vag0FN8bSHwLLSS4n+AF1oh7wWJ7mOwS+U2ESHYI/6g581gvAegEwKD+glcnKvdkzz4l6k1veQ1R
PleCevQFLELXJ/ZUMDAUaPYsC/wV2MlsHu0yJC5gRzHwzNo8r2ub5hWX77ZaLwS1V+1wJuVIkho0
/zcm9ORaPQLR8lLuPvJkYrN9G+y8h9kaNrea6xTDJU5nOqbYmUl+FV3P/voUQBxrNw9S6pS3Yp6b
5y6PnM2hCzfIcYwOxqhA6cQ3A3r+sC8bk0yafSxd8VyoLKrE49KXB541Q+t371vt+ng3C0v9jWEW
KHUtzbv0lHQJ02I9a+6+y737eSx6wbzFwa2baMRMkGYAdutF6JK4rqCgYkq3uLtSORRi0BST+q5e
QHmfcGi5ADiDfkHrREozVfHvkGTXoYIjd0TFZ6umecimZ+cdCuyBYDrsS3T9URXR+9XxxkWyBdie
OIilMbxT+S++NRs4uLdke4ETNINs/hRzTp5gsrT0JDfhZj0C9swM6hAauSw3c3KPgTuBdhTKP5aO
ENlzhJqUI4pr3EGctCTtiM3aGxOIt5ymyrx3InwQM7HPo/PYojDLUqobXpfimxbYXad3bmTOm6a7
1xTahGp6tcc4e6kk5kIW//EKucnmeqe1OFEUhxgV3FWqNKXGiuaVfDIkuG6zeoji6rNCSpFdTM0L
yfy0PlPMocmJm+/VWI3gPrsEefmvyP/UQQ2oyDVThG9Iu2ItbF9XhFzMq6EzbIWG22PITj/09kXf
vKpgMw5sxl9SHJPYNA3FYmdaxwA3BvQbl1EhXJokNIVtiV4lpeQq8IVIy7HfzlHYtMRc6sqZ6QVQ
ba1K2AOoPI3areAid+YTank7uv7fiD0w9xsh0hgVKZMr1wTPqdbc5Db/haCMRyp+D7WiZHrFtMtx
vZ6Bj9iE/G7QoKlY3AalHog/czRPGVUPd5b2GMwyoC2RTi7SVsZZQn9Sbrxv004EyBe9FCkI9Omd
Ss39PeMlZ+GST+GosVBy5WHlhLk02KOBGaS/Xjb/hjR4kJ9Ro7eDgjSx55lWZv+uWwRAC4ExOzP/
uRBOmIQGhYA8aFIGsOhm3E0bmZBw3lJrhEDPhgV4BQFXy/2qY7KS3t7faUUGw2FKlDM5RAPFohl/
GKj7G+tYF1IAm55tbAysf+wKBUkjtn+HVSN+Hsi8PK3sbsX51dOw8rRvfcUIxkC8TDMVnd8ERo1e
PAstC6pdsrxuchIrRscIi+59QHwPFRxDijcjxiUTqnojdk69ykQP55jHUL1bp0B814kCucYALC+c
B8Kg6a4YinS9j1RNcJVzM+WJeyNhqwHm8Foeu3HJhFChefVq2Tc9oaYeMFTKvXwVZS62/x5qnrQp
EV4sCH7bzty+bnLdI89ofNPUaxJ3mSsGiZgy43MmnZNGvRsN2Fv1TMZOXmRFiMjN+NA6HpAdP5As
2fS8OMGyZvw3GjC8VaCjOyG7ISlhd3zIBsUUVxV7gjVw1A8CFNT5BFsKVE7hdVkNr4Tb+S+qrC1x
kKQDbmc6wUkTVdDpEO4Kz8wKZTxp59NLHI7XGQf++AcwQ4Nd6wyxd/sEg+DFwviRmMrKZCSiByo2
CvcpnjN+grmfhdTnWCTEAa3zfQM5qS9N6P34qSzHImejS6XBW6D7RGuZkszwZXvp9l3LjQqiMRWf
n6QwNwj6a1GwaiEDeBt1EYih0W2jZNqSbZhEZwdS1dG6hm7VMsPlL/melZS5JfujumBRePZ3u3c1
HIRWeGpgBWcqmAayINYAwmDP2TLrj3LZFJulSLZIdf1SkPFL7utci9LQi0t/Rn4RT/imRD8rVNXZ
1cZEQV4R5gtAkbINQxPeWJfR8ZZooxQWbrK1zg1bxCFXnnQArRSfpk/58ZeG1AfskVX3HtlGXzCl
OHfGnhnvjj5vYoODrYSCnmFkcfqObUMaFz4myzNu917429JAtm++s9LDeX9O7dseSSzy11xk/0OC
lDBtrS7dpjtec5k2gDmHAo3waJ9H/QLhwEzIslp3lL7U+loiJVYDYARNXsGeo3kiuj0OYp5z7BkW
ar8bYY/Mi6aBQIbmoUcrBNginqfeoUbN+3FDoALJDI5sR2GOPu/UWTObvhrOqqNC571ldppyV9XU
H/x2qvuNvDCL9XC7OO/zbEOevLNSAi5SZvm6TJ4QW/G30BUvi87oqBIk9C55BHjB7PGttfGDMrI4
mwfH8MYVmPYPFai5fB2MBJGS0h9XaNIY3c0Af0fO33KAY3HQ7WcLKBO/m+K9N7dFRlXpizZkRcL1
Q98HFqRHVavgpX97Rz6l50jnl4svrCvx7kyJpuxqZLPYWn0weXEbWLm56QsUx82M3l7UktF56eei
ffcCSCOQ81J4zfCzb4dRUrw7zyR4QYu2gGIibzA9lYyFKTU+xW5kyOM//l7mU17/QXZGlPt43XjC
u+/U0D4EOodDAgciyafVedU9LQXWTqDs3xQmWv0Vy/OOugh6cpFXr6GxCp90SIH011M8gJUDOGCd
OeUbeGa89CNTwdIk/kfSbtjQG+PZXIuEIK4wzzSSx5+4TevGBIy3ZSyGGkNrtoI6CjyiDpeFNrht
u9uHC1Xvv3pYro8mtxxlOFXABdWcST5z9sK8wE949kfJRh4D5FcGi384oUAwzF8WTVGkuPU+JSfy
fR+1VAw6tigbhuHClnvLVEH/jYzWi8JSssDEN8RQpngzuPyC/zyBOhHdP6lc/jIv+/tEmn2S/kOe
3uGtsIVyjDOg6PNXauAnYdlkerHc9gvlE1bYALRgIhbGyjXfNhJ2OKWFdz13m99k+9K9ebS8mSaQ
XpfPzdPBpJCAIQJbHbCvz4rf2HvhbF3dgzJct07R3fRHGSbrkBNJ5SO+6luti2fAfjVUOsDCI024
lT1kfVjLK7VIKhYw0czKKKtBwxMaSCXAbOhzWvVhTOTygdsXLb+mam9LcYuRH934gRIivVJ5m+5V
NhidIt75JmUjcZ11iguwNDhDGDqKhz/d46amvb3arJwmMF549lHMZ/Zdk7kthEr/BIb6WNajSChz
rMknQNjSDrCTBZqNnk/34DSb5hQzUng/Xy52GNaXBfTGbSMIWqZ96ZtoLVlF6CJxv57abWWqfITs
s+JGh/bFFB0yHP6EYFqXOZhxH5WFtwQG4xWQwUG5mHHOXagOByNmg2pbH+25S4gvmDVcb5eBoqGE
dtGJKbNLcpgBriAxH2tnSJOQxG9HWDUmsZrzj56CPFK1PNVCYf9ill/PEaPL0TpeOvhMNS4cFq1d
M/wGtYjvqVlrLkRwp8Joa9NrI9XwUSyRbNn+iquE+UgLTyWEZy2bL22NRSwquBc2TTThSFx/qnCa
km9KF8I3nClhPaZCBWQclaslYTi9swFKypbDqTXIR/o2Dr0f54QMiDVV7lk+3/bHLkOm37FjZoZj
EQ3JaARuIu1F1jGc95Uk9P9A6sKRzZZ3Ejoz4WUoH7r9/LMOh02QKiaZr0C9oyD83v0ClAvDTZbT
vIZeh1W2WwbsxRXc5rkcptY09/tI/uS0hhjWMjNuh6B1GT5KPza4UxIedPxDPmN2qBOGv9JENDFc
BwEO4465sCtD+nIC5wcaqG1DHazMaFz5KD981lGt+afu+DHrtKppU1XsCl7hkrJGrzl4R2JrSFYx
ZCfSkFNiPks+coc9DlQeEHjj+bVTcgGaFAcG8FJx3DM5RyX55oM4gH+JqIRNK0kNo7KPyMkQqPEj
inSQs0ATpGOry9iOy30YV5M3w7nq3wnL6b6/M7IqfblH+feFpWt+8g9c85AeyStXN0+qey9O/4+w
NU64tiaixr/8Nn/5Osd6QGeanpv9tNYRkHuboM5SWhWTeA4wyaEsQC6uY6aP+iIJ3KqpCP+BbQR4
Tos0xyUWSlZ94MfFy1WNYaEvYUwEwJXQCxqDPi84MFdwz+7/sS0Cffy9LX4xWMyDtIqKGMU2kLbb
1HhlgoPXpaDCrlAQgeu91DJDc557qMNZ9bzdRUKYjHrNEVjd6eatJISnDZHTYGqG7AAgJbqz88RI
JRVr8ZkX4dQtp6ZmJn9933S19KHPwSTUfW6AfE0o03HFYRNJDUqlsT9Wg93AzILBhEjni0lCa5l6
eucFFBwPrsMOFWpA104DAwQp0ry3J95Q7Z3unXstJzf/dbZfsu38uHc4Am2D/x7c/UsUGlSSvRX7
DjfTvNYSYqoMt9spYmXR04lnAru5IxMkxe2IT5YU0jjR1Lc4t+G20617tX4opE2zrw24UzePrYgG
Etkrx10Jf+tR8TlGOPZkpNWavuwXhrHsVzxxKnbVemkAuF8MYqEMNQvipTPaFkmFzLFCJGikagqN
L4XbWyI5d7CICPO8B9zCudnUF7N2K4TaxgkrKm/kwFGKqutOJAkQPCY0fS1UevXr87yRS5N8JdJ6
bO3h/7BVaVdhblsrQlnj3Pm1fBCrqvpu3SydElDvv8fwsIfPvzz+mGgDqLb/JD9cxs516YiEAyMP
hpMHjTO0loj5N7qi2n533ppUr2v3qexIryxuBcFWregFM+AxDIPkJA3arZYXHe1pKnVBqGKKCXcK
3lEFedCDlXPsgVZ3UlaasRXkCRlhEo6aOiAU78DbeHV9sOvHGxAJCl2dLoo1U8T1m2lr+4dr0Bmd
H87YCtRwJr/zC12zRXnvYm9gkoUzsqG9JPb9gyQ39X3hkn62Z1luZbid43hv08LM3bnvZobkrWYa
AtuY9d0VeTnTK1CkwMNNdEgbsNuggppeWIU4x7HD3aIydG8k17NTUmRpIDymQqGyroCMss969Njr
nRQr9dE37NiMMkYgWbvSpn71wORvJnqdjwfXXV4szLC6g4HcXRjTKvxq1X4mn/fnx+vIs0PvhZ3V
TZa+FnRINavzPvjFF2t0vMJBVjrhIWHADnAq2wgOoG0a3zvI2YcY4H0+5AItVZG8da0hRfE0IdRz
IaZNc2QbubgP4U2yScJbQuiKcC2X2+qUkyCO4wa1qS8EiJnrXKYMdb5In2tsEto4Y4f9CJ3KHXCj
szy08SynDp863NFwAyg0AVfG5xUXa9kHsi7dVk68m0sfZSdgZcJ9Zps4swonUGlDzuj+rehBjAH5
MJbNdKXmwlIzH2TOqO5yqV5Qiea0Yh8Lbg2ubnaQ3+2T/zuBksUcTfP/LUcuseAwTzdcKtknwIsV
9oE6nbL5+Tl+ylqEG5bL0B4+biM14uxE3giRONnM5mb+P6VNl02rk+rCDeSYlpD7wKRnwTV+073B
6YGOLKeFkKX4aERi/am/aHX4JuzHQafsR7CONxFkS1L5g1J5hDjJHBaQEo4FQDdKbc+DeAFfofJX
zwHzdLFBSq0jXdHNKH90PLMfqwH+igy8jCwqqd8B0uM98jjUQrtaL5Hwf2Y+ngQCD2HpOiLbi7CE
x+qB2GOXxrM+ZJAf6hyac6E5UAzKvM0PXb8TFrLwKALj61fCMX0/4GUXhbktKPuiJ0mROhaDR3ub
Pd6xmSb4G/4/rv4tcBAOOSzx9B3HK33Id5BRyQIrsNe4yhpwb+DwrMFOpjtRXiGEskRmi99yRDLi
C2eIz+FYliWF4IuQ7CIRsSaeqdRfTlPpN7od3p8MeB83CC7fYgrDc9TYLmnWdjMLgWkTVbsXNQPe
p00n+sTgE1HQ3VXQLtJYyel3UDMQkmvQXiFn+18oEueoxYW24SDkrpCc0ps8Y0kSdHT3nGOuPV8O
IrYJWsiowJK4n2TN0vyAFhl+7aS6kxqS7wtWX1EMU6Jr8dsmY7ZBgO0lo95eeSZPom3XCMppEdtO
fnxXJa6jK3ww+c/pWzG+YXZn4twAKIXAUhpZMPSNKQMQr8s+PGySJDwfeBjchUhllEl/GwB9ttZj
hXLd0whfyHDEV8cW3w37oabsrR6z1N53GxGtYQnc4Qb/zzsgJgGhtRCPjZV/8FkJVUBjGk2nFUDg
+jP7Sf1muS/broSI5QezPfM2vC3N7LHLJVOS641wcNnDXoLN4U1/D5/b2YMMK9FlCLyad3Ft0AtL
wwrSUqUsFgd6hMuGAUDusNO6KcG/waPYD0RGqlOwfdVNBCB/jkxAMVkkFZFPiTaHPrP89L/0DGFf
/YoGO3WOG3soNhdbn/hyCgLTHdErg8sHgl7oi20/Fp6XtuzPnFgJt0NyDA86h5cHL/blSSr5/PkP
OpCFum/xL52kh6RwAmMfeCQDHlAJ3sTklbq1u6+e8+rfsm7LpdPY9JyGMnRYc0TVQ6K3t6tVv2Pm
Yc61wn1FLKt25ovELQF0wJJCXjAFkf2DuMhVNGO1JmRiTsKrGfITLk/1O20prwn3Ipwc9KW8l8HR
LxBs3ozk5vAinOEPR9DQmGOMuuFXGC+PyaALmcbJMewnQWpr8e4MldzaHE4QVytDZzlNH4E6cCM2
GWm5CD5iq4OYIMzlVyoFTtcMCbtwED2KliWa8sFHnaH0yNJtRBbeigbAp3CZV/nDiMsSH5XXz96Q
kGGwtExHDoMKL0yTrzvo0Lmud+TVH8xWyuGDsxB5LxMZFfD0TmHekmth/AERmbwZ6pTw1AUp+PEl
FXDGWps0Be8vdgSuzi9gN5ZenWADdFPqUucaNtH8ZXCQX85p6lDg6Fdmk2rsk74xP2C62zs9gQTC
vXIYK0a4/bvR6zzkFkmsTUDUjmiBMsIimWBF+O1gk0nOJyE0mAZanB/JrP1L6C7hT4jW+uitky6C
sWCJ1xwXaEG4mDU/OZ7nxnDus9KJm3NJg3MJPPiV/YGGrphKs/xGMOGj9nLwlWJG/UgkKVKc+UNu
0aztt+dJWYITytQQ/14Ishyy+vKRwDe2gNeOH6+bMlLxmXkxnwsIWbmv9e8Tw2ezo+odHf/x301M
6wcCEczF/74CHwSfN4XzB/6YRvDCHlFME8rvvMecr7QJE5QwvFEQWm+mtHQc5Lny2300muHGP7W4
7e2y+nhHLaIbpXq1oUhXCezfda4K1qo8fZElxWGPeEfwVgzbfa+1wViyc99Pho35USLckKN0Ck5Z
vKw792lKr0pqGb0wKPM0MzRt2LyMN7Bdmxn6Kz3kCCT9FM0ay8TgXUJkc7eBVLTcvWeZ5p/xlFRh
5CqWqSVV6ty94HxBiP0FFneCYOuZ9BZwnSsl1mlfpSI7IFFivgehQQ0senzCZcqjebN8mdvpXMGU
CZ8lbRfb/z3LmkiqxwKLTeik02pED9UWDdSKBBT0bvE4n6O2k189FWhlk+PLsncYpaaoFFe3w0ut
ygMxhhz0gNbpliKrBk73UG2JmoVctoAuqdky8ECKlnEjYLaMY0wogpq2G5fu1CIFBNsDs+IKKP70
jE6ojLNBebpQfQUtxI16opro0+wV8Z1EkWiLu6FXanv6mGqbGuW3kiaHDYtiDEBgPTuqGwYIiQU6
q5KnNpZNvn3gm8n6ACwiVtizxgTd9Gk9Jhb1ogErDUTxpza39jW48DTcQG708GdcLSNQVcBmG89f
GsL53duWzYIS+JSnnlI3YOENuROa+YUAz4I3REZl74KUm5b5wA+9c+01CcYnZFvRueel8eNdKDXA
NB2ix7teL9TVdNQmlHf/T8VRSOEtc3lvOA0GA21CvOIq5qkyq2vlXiUOT73iYfadXoJV5b2+VSue
9sLrmTDD9OJgBLYE7FM9hDO9hOyLTzcp3XVfAkc17i5mdoUJqd7BVvqUEvvAw0Fr1urWRL7KqEzp
BgVJ0mJl+aUk+NvBDbRqawrdS/En0KJX4S9EayiibYr+gt2thHxyPpNcsfuSp5MR7FktN0KH5xy0
KNN+5y3Ki1TOAEgotHU0nqNP+P15A2aRtH06+voX3/lx+xtpVFsiqr5UCdJki9WzDQqGn/TaW9/C
vx1NVirnHLvyplQVgQ685MBdnYEIzps+1CWGtf3SNVrfNNluqJj0fB3fi6MbhTY/j+S3pmTkSDUA
VLYRFjl75B7nRq6TUg9AkNUA8+GA1kpnFlAzXpF6d+9SDYZn8EzxhnjFaKtgpr9SQRN9jFNZvklm
2d2KQVUl9onPL6XmVmdGhtDoNEVM8Dcd1FNtoOwNzfYnxF800QcYli1EsTpXzMr02LHWdu4ZLNwL
UONB2lUwHAiIiuy3gKalIw6KHXYIijrLqeHeXtHh2WcVp+9LzAWbelU6riX71wnLB8aZdxS7xYLf
GHsRr0rgnTRzymMc/R8eYzArTUqZpG0tvR1h5Epy3qyU+hG1JE5JX9MJXAh+ppfj4XU15aezLsOt
k55WcA0SwjzGXbd0+W5Gy/diZXXLbZxIS/CxVoyOzz6bC0+QEvwxFKpPUCfcEneHKB96p1UXKEEx
Nzd6bD+wxXqdPfCQM1XGfVkyKjFEBdzLcrtUOEJ3ExZAc6dLhoAMUUUgfb5cQ2t/gYezwcpIWYZq
gu1heoJccHCCq/AR9aRzIdyWVfVMGzSZJLlIPWK4HQDWRWxwBycGtyWWAJZAWV/F4txm3lIITe+w
oae8Y0Hd2il/fe4Iai/AlNa4JxnX+KxNx4IsNy3VdmLYuXH3oj7Ez6LY+O1tTtFJaUKuZb9oD2cI
u/XtaTjVboaHK+4vxZMF0X5w6rALTeuLkHdUyMaYz9LDZ2OEeAEqedw+R7biKdcNKEM1RTKuP+4z
9lnfyBIhguCgyKZZ8PhEBiqInsq5LtSCT75dM6SUI3J/igH4ZtVIlxyI+87x1MeBZF8A5CgTtjJz
Jcflz+TbVqUascbcBa7w8dciKMG0caJEaSgb49rcK4oQlFYOdwaeX7T4cUtf7stXR6flOf0bicd/
aD90tVVT/CbG0PVIDLyvTEnUpU3q6SNPxfVDfmJaesqGPF+23Rl1BUN+l+7cHbTXT/TzJMegwyQx
mZEPPCkuJi+vwehxSeV2k5JcknulRDX/kNpgpX7oWuzcX8PgzAn0eID5gxviCQzHjhqQwR77c1HS
8z+ZlLGW9SPnNv7FHteb9y/n3bduKoeLbHz0gZOmImxfFbEBAGnIwWp2jhHtTQx8gX+nI2AUIiBk
/qTAWT4/JyTENOTz50YRC8JdLjJDpsNwScDk2FZH4l8pZUVofsvnMGNsGkEeGQrtH997q7+KN9yY
wfGinoHvYjDKZGlv/YkwQDjVEYcJceDC1wdvuP5xVmIWsRtfgw78lRUvwJjz6Sog5AMzvAAOd2G4
gLHaRXU9bHsN7c8fSicmbqC9WQTPHDb4lsrNjr4odDhFnZmphi+lkvg17/ExM5wFKzMyhioAMgbX
pIDTS66gjl/34cOBoe6qHlhiKzGhQmRnQFchSAGWef6ep+/91IACX4ttmWXI3Loa+5pN3DTYbbtj
iJmtR08gyVJdo9e5E02buvB3Uct+bg9T1l5vibWP5nYDb3c7KzuPlL4h5ruDKFaSaMOkaEIMpZP0
wG9bxZlkpLAlXQ3jFNybXbGl1Io8WlWYwJ1mm8Sta+GnSp2JDabD3ce/UVa89xsb2IL2I3TlE+5C
lCHYRuhLzJCzTPKjybvvJJsoQwS0B6gM6peWwL35w055scePwulw1EdNRjwLXHIFA8ETKYLCbtUv
CrArgYTi+lH+5AS4o2fh47w9Q69d/LgtHNeqq+enHUQf77Fc20MrqrXCtglv10XvxdLvfXdjEiKA
VMJxiP2MknjVvP2U5vtw8cy4ddKuwvx2b6xXJ8gRtIMVlp7NzsFLgNxs1UufehIGAaXgyjy34kuT
2vPUdKketuxRZ668LIONExEePvrbwNQ3OL5WlD3SAXK06xdujZYrCVCEsz1JEYZyqJavHNR4dfQf
oSTXcG1M0MVuQf/s4+jeo6DcVot0k4mfDhd47H+fcVJyZa8F3f9rRyGbk5Jvi2qeWFsTxpRH9mrl
ESs0OyD9hqjxLwOKj/RUPP7x71GzlYP9rdwQI78LLyb4vCxiRv7QE0Dx4Ly4xOkFoaPY3LwUXyiK
uD6ZcvpTJq51gScOwRjERNS1vSEil9gRuyxA9f0ce2P4kvsl8a4NflrKynGNCla8Ey4YdO6FzO5O
H6I7YSO0nOOz5EFUwFyf86iTtzKs1lDTq/8A2GgneXKIGmQtaEGsjiexqid2GmYjKkWBetd1Gob6
gZOs8pnc84yvaaj1DKeQIVKyznaIWAzNtU691nWhoXi9hrU2pNBx6WE98kpZFoFP7cCjumoW0hDR
/54yPPTl+Gpg1/YIhEJlTlvncs4d7Es750Ek+EDG2MbJC9k/ORA5YIkkzUQJsDI8c7+30J+odg/q
AIw1JsyVDnTcFZ9yaLdzIaKOxMunXxk+NMP0wDrbHkIgxAEvU14Ps09driniI6yL+q4wHhv2aK/9
uyrn9AnMyaib8F6M7l3EbWGX5hG8vWEMt//aaoi0czkqpFcNZKciOnOuHeG8j44+C8bAtOZfBFEB
pzRT6xSdQku+TgFHoVzw/p2LpdS7Q+dUPZlKCYYRKHtWcPInfR/xmUyq+LviIQtbudSJq+DJ1ycb
5oSRL9f3CE7zMbG1tE+mR+DACk9X6KTfyrKh9XLWlBBNaPNqRVWjG8O10feSixHzZRK+G7AXeFGK
FMOCGhqM2uPa3spgR9+B8fFrWo0kQrF7rqImgmSdzO00F4cy+jFPWllFU40NNnQp2vMwCuovNeRx
Ask66yjdCsM6/h0s1wZmU4LtZpxC38P1bGskXz77eO/grJ2/hJpW+/28YKjsDbS8lUC3lw7lHyYJ
zzNao73xPL7o9Bk+aMo9ss17esuNb3yuB2/0F8FCnH5It5b0bcoRSxnEi0c4Tw3gRcJ6XcvlyPlE
IGhcelE1rqsvMMHcqBvhn2F0hrcbwJ4iQYiQyq70jSMBOIWtpzij9vBzDAZVbrm2wjBCB5g7yQ2X
G/SCplYQNON7OseYqOdTIcfOajcmTMzoYa0KkrJVAX7WCCofo4cRUpMiQrMFWQ7ZapjXJ5vmiU6X
yMrlLB04ppgbcjqxRocxd4QWfU7tCAigROzbMMdEWc18I6+59mLoCy6WR7iLBuJSEaI1oUUYxGaR
ux+XS0fIZBuN4ts5cx3w2n+hcswrQGH36A1hLXy3S8Zy+qcQKZenEucd47oViy1y6l4DPxQP0TY9
Kb5d3toXaIZAdCNheMJrC9K6dTTWVglQ0KXHyiGEKvKD0Ml4HLno8fof7pf7L6Ea4K2F913yv67N
Ce7YwakcWp07Ln699lJ6jAY8FfSgAqUkNH/jfTaLHf/M8LaMJisJZiJFL9t6CBhuQz11cotdDaEL
9sfRA3uZbN3ofSKvA7Y9yNtTVLRTkAQbq2sK5QNCiaVb5PK8Wuq6j81mWlCuDaiE86BFr02lINaW
FsIFigdWK+NcI1uHTjYs2RyP5vppLkfhigLwhjLdOtAnQhNo2caCeMa3AovfH/Cb/vBl7kF8fNMT
vtoFVS4TwNb4d/mWPFY9uh+BZ36pkqkkr4TmUHl+UXN34SefRs43QY8yogvfUbFGXxrRxxETtmpT
saKwYYO50WFGffU1waGsNWDlECaJMYZGwRzu0M9NN5edV4UbUWXZU7RxgBy5A0OqvGYEp2IKeqmW
mrtxulazUgmm5xlahrRpV4Adft1KRxRqrNiF0rBOAYONEaGA4UTJD3XbmT+Vzq7dn/ZhVHmzJ27h
9Y628DvjX8t5TnOhqbeMNN+SmFQayPGG1Xs/5uobyU3yuVXMZGMWfs/xqf/LqnEeUZUxgG15rqY5
MV2WQukTjk7iee+1Wf51GkQcvZm1z8ECRrkhnp4FwrRLtWlwQJ4V2W8D+Rn1CwpvL7yElNzah9qJ
GQmATxHvlXJVeHYV756/GgygvCzwfVfX8U9w1uUwpF3WFf+RtwPZix6C0DYgpqmlYIUOc18Afiiy
dPM8DwWPpHdEqlQ2ldA6VihevHQxDifKHhfqyfXFqaT5ZnUVeyV3BkVJUy/1Yg5yByEDiLkoTQgc
6lYIEGwof3mdnFgRu+SvPBCt8V2KibqN7NJ2Hym98QoE91R2MTG/nkiFJXbCCHoThQpF9GRLnGv/
nprLqurCeYhN+Fa+fa/YqKnpDX7eXMER65WHeq21sALGVEgthf0E1ws//bK1FOxPEaTGsNtJkewi
J//O/lvt+dIrCU3l874iYfkqT7sqi27wC09f6plmXR2COYlY10hu2XcM5gchnseT2+fDuxPZAqac
uMrazVh8mp0fs5iqtetlPzEf6OzUSTH2h8tckoQCBDiDOCoF5laebCR3kTOvRwFb9WYqmDIdsT59
M0IerIHvvw/BeyKG6hVyj7Jjh1ofEcefM3yw0klOHsje1qOOlMynwq9CxXt7vpOhhtleceRM/e46
P0gamQHwQsPYn6Dl94NLtB2Bpw4oZes+qGInrQbL/h/qSEfJzZdFLFTquRwV1uFKUAo9O+MmpvWP
QhwADPrENW4TFKuv3Nc8Mmvaru3aTnXY8ZqA3H/LaIYsy4v/8hJ7leRZoI6EVu3h+hnzsVHHraoC
r4q/Fqv/4pOQDEl6nYdEZLFvfJ0ekiVLOjGEj04lGmRZ0h1I9iPccVrxsxYjDak26QGwrLDxVtMH
/z5UNg5SeS0j8SU99eO0cW+We0nu8fG56EgU9JiJFK/9J1VPNHAU7sgQB7/e7bLmTD8wRtRfE+rE
qHCBeSULiUBRon7gCFg6HcAsMNmLfrbNQykTgYwTpoL7srpDvNgKGtWWisC1Fgpd02x/QfkXjQ6Z
oMvlq7/BmbkdqL/YIqNKn5tSEILmfx7YlGKutUZ3pk3+xuDTOoWRs420eevrVgeuChWQITRsxgm5
7beQS0ixi6tqM5dZqAVk5g2f0lEo1BD66uyjSEtdiBe0qCzqvcBUKH3xfcYdn6pPPgSlvhBiGsZ3
tdx0aigm1R+PedmW5HueXo/TZPuKutJezRHP95z2q4fQDfiwafPfZ2x6tMrQKuR7JwFmyEFTJqc+
XYsvN3ZtbuJOwuYHM99aEF6KThZWrdu3VCW/lnSVtQYT4xLPD9g0ZQFEqwAhNL9wPhZPC63o8TB/
THDG8UCHWA1TSxGC/H3PuIQGEDj7APxbKHBWi0tZ8OFPzY62+OX2FwgVYcaDMRdEGfE8sqT0exqj
H7eGcCczScxSgx/C3ToPA4k7Sl+7z9ISVaAgta8sMzRJqwXiyTfInvaf1S/l4gWKYWk+t6GaqxUQ
hvQ5kPDQPNcsTlpl5rejx7HYFRzLUvWHPIA2ztUPJSC4iPyXUDvp0HefW82zVykNxAVSWtzohOrf
YUvgDDKgX6uomQex9JQCutA1eNhDsBKclCxzbSKriuI16XnoYmaSEUQyhWDIK4wWHdkadBZRrrMB
4qqNH1vWneWKlMCK9JMTkbOQt6rBzEuWHbIFI0bnBouj0sbN7gM7GW65QM1pC0k5ii97gcIcuaVN
JsgZe8nzCGybBoDoE2Dbg0esMJB4xIzLYw+H5RJgRTbXeTLj21g9YIKbxVSlHIVhgwTmTJQF7MUJ
7gD2uTWArqb97AafqNcVjFYuhGB+bnzbUKCcJ3re8OkhdadXHHD9xJ4J4PI8nJELgQx+51yzq9YC
MK2LLqB44Zzf/H5CxOy25fidz8v4sevS9Zvdmhg2nMM+duN6apGwNadKZaYwXC3W4wgWUdDeKxYP
dd1WtnFmHdKeytRcnck4hk8/9+R6EeO4gj4eYXGJvjcms2N1R9lN5wJ2kDkJAC+BAvoc4faJuOhG
yeiTM4t2GENp/WrRlP6HTj1gNIokz7mC/HBRCHOXMU6CltLnut/0IX9IN2v0e546s8PtplCGFSOe
Shr+Slgy2XxMWQBiG3lqlrahWppnHkd8Umw+nnl3mINXKa1lIa6b/Ec7OytkGRv25YZmEoJ+q6jL
48BXTrzD1Ct1rfWZacBcd3f8xwu+80ZI0tnjzy1v+WfmGlrkXSQkVKSMjiarjhEFTBAHSw+weki2
81boTejZ2NmNq/bvjgwX7UyvMspc0eRGrv6XzitZ3zGHsgxUit9t0Az8H1z+log67m9081F4D9/C
fsdaaODkLbc8cJUtUC4Q4j4jCey8y9aryP9Qyzsk0nRNA8POSlVfnlbBepAKQ2hA7jf4SYpCRWXJ
ttlP1JJfaWpfltBB6tA6mxAQ/UTh9M83m7jgE31jf1zIOMBv/v4aXhdZXr8FOCvBYJ9sEXRAzvUE
MEaRshav9C+FatiP7Fc0RuGiZwro8kCei8BwPmaJ9G6XlGZZ0TfCqErp8H51X/mU5/MF5NP7yiAP
cRTrKrHMAvcB7PW0QF6dwdUH4ORaGNwQeVNhjFgi1rVE86XzPwljj3Es1LLKpjoxDivMmnBeHs62
EhPc0dtLSyt/QdPucMIx1vOLW7v+gOlByXrb9krqo4P2nSUSAJVq0zRDUc2t4WAXfdatu2HKhgIw
7UcKuxl5lbEfN6ReDrDNeoKVOCbhit/qLZU+S01zXaeaxPNA3+P0v5BmNgZdUG3vERLh5r1UoORD
7HvJ4ntt/u+DnpdYC9lnGJFCdqyRUN4zzqHOcrur8nwIQok1fwxR9ehHSWUogYvUrPRyIEWRV5IQ
BzC3Q+Q2o94jE7QmfRPFEnTweYi7dwOlmIbAOmWAARu3CIQxjY+lfEmTiGow2rPNE4WyvNt9YnuV
UhiW56WlYa9rSOAdOtnbXD+UuMsV1IaGAzOwO79iyGmjCapR75ltNm7JqTwiP3WeCgnnVXYLdCKo
Dka0ItKzLR6dMFkwvWGtC52mpWehn4oJsNYF2kwnu135AjW4cnDs7Y58yV36AWXafES4Tb3yWKgS
MkmzUIrVt+cQcEqjV28PbdD43Z4wSbJqRVi4en5fiRN4o2J+McNxEjZpQzD5VPbY1uIwmPdDxTIz
tI7RUQnFk7u4u2uqB9VWPwOVaPV+VoZqkpo2jD5YZIIjkEYjkozHB0ea6uKputY++Lie6fTTRlmy
mZyGG8laUecj4rjb8T1DyqIPvs5uHS6sczOjXVKXUSevdFqyHvRwLC/+AGh5DRH2aX3pp69Yk/n7
Lg7hI4+HYZOaFPGnwQvl8xXcHltM+du6+hOj9Fn3OIpTcE+wMm5axlTmzQUzWQ2MwTF2aXVwqq9T
G9obfUVIPqaIdkeZuONLgKsrEgAoVmlLm5aeUO2pzo3Few1CXoQ/SUl620tzg/L25/KkG2FX7HYZ
pSi/Ik1WqjIlz6YS2WTwcD3AxtjKTyVkeCaQS5yBZjuGgLTfXC8RY68jrA3QEf/tGwLOU1hqeJdt
n1gCS30L1DUvHICSe8qkSn/h6A9AiW5PnVahbGOlj0iFTEzfCAlaL5BZLyXEeRwv6feKFTPnLsUI
cLktoBaYWIigEzWBte209JdicP0hwrz7j5c95wTEjGT+ivPRzAH6UD3xT0baVoBdHpIEoNRN8eCw
GV3EbnLvzjQLD21p3sieuG10j/cYbsmzVxVXoHqO7Kir0dZW1stng7Fqz6cWoxLH225qYLzzhy63
vEAR7M0USoG+lOxzs1L6emZKcS1g8YNLhEZdEWcKnft+yDC1yiw66C7WeLUk1tw+3kpeDSgagWj8
0m+uwWgbmu6yZPnrKUGGA0Z7Nl76JdMtZetFe+zrckRNrTQUUYZeurw61yGrZWowy4nTHJzyIxvq
OTha1jhfRzu3336C49+gUoy35fH4pNbu7SV1TCWxnIdYhSil9k/6wckpqvhWwTAu5FoFLrVJxlAO
i5tMvUGwYy8bHt+T+I8Ufwllu6QUReeFVgMq9MGJWrrQ1HLYFZyeogudvCLDSmTe8p9IK+A9w0h2
e3HS0ri+PXoA3k/qWJn4Jouu815GPrtz4OgyI75q6owjiH0h4x4h4/CcRHLMas8eiC1kZh6gKqe+
0OxjU8dTcH31Gus366oJ+y+xJsR/P0wmcJxZ+ijh2TPduE1ztCDbTup+qt+H5OWy1fQ11ekpW0tm
gjYadvmj1OvEhR2c952+MkBDdNi1tI9jdMxvNg4tYg4Oqk+smzs3R4MJvqzqCro2p4UjxZr5xNsy
1VMnixETih79YR1CcGF+54YIgE9uJV8RJd6NWIe9lqP9jPHfCwphJMc5yZWpY8W9XEmTyE+Tmw3o
Imtlxylw1lcs1wM31QvNUwGpiPAV9ntVlBJ3Qwad0RyEMtJA3kvrm0b35WEtAEHMeJyeVc1AjJv7
FS1GTx8kCtzcKmerc2DMFxUIRdj6epykFWcaAJ6KniVi2ewMUR6lvsXK/o1ZXTYKx/aOCJdAxivm
yv/gBGkP2Ey8WogTiWEAAfVWDFNeJ5aZ3ISgknI4K0nMZdqUNcGxSB7/Zrr/rzuSE5c6nvXQ6RFI
JjB9Lhq7Fd2Vm/Ky7trU0NbNA8f8tYDpUJxEDmTAMoFkHmzuLf1BRqffFAlZV7bcePeNgidcHUyF
7v9CYZtVQI404J40E6jfDghKZTRvvOtPeMNLpCcGxDMmKi3UCej4+gga4pgnRh/WlmbYQ9eQ4UQA
TdtQk8cJqsZ/OdPdNV3YtBcq6q9pP+3Cg6QoET078sOmzgqRkG1zRUKPomNGNAoAiQcWDJNMbTOV
3HXvoMfJ5s/JEKhrp0VQrSq/4NDdaSswQoWUg5xvFdnWKKr8hZ+hZCbl8u0vpMxSb/wiFQ1T2lgE
awheZDxDSYhWYwYc2EPujWeqXiOG+jKTqElzwKTJX+dzMIWg33Q+GJaxhud08PiJi2tUOHQCdBDo
MdL1VvVeSxuB+2HUKkGQ7bHaFZTMZqrgdYasxEK0FcP7pH2clCDGGusqsmIIHF+AXYe4VgeYQFso
X3eKHwcoRzaPbNCYd56kJ/aTUldqKowoxPj3/MTJdUx18Xk0BvbtE8xFb2ERaqMV6iklubuZlu9S
lF2dQAvDtRC8MJBchwDe+oY2DF+yRH8KvS4BHvA5fuBdaxvY8Yl4tgdslGy/qPwpOjCSfh5Vi3Tr
5fEqiQwrIOa/b7AdWaclFdaLmRM7/UBsm2MmVLp8CkFFaU5JqHAbA9Rxh7bJqN0jrscqMZseCHDH
8RD5f2qv73+0zyPZzzcfw/W7sqtiGQK6d2iYxwu0lpgntZ4yYZphMmAxdF2UyS4wt0nSRZUyNW11
Ua4903PckMX7cACOzcNe0jqsZT8tUN/RT3VSGk8k4gZJdG+hg4gDn/hwZdXmZsn4iFXsK2q24A5D
1GZQx2OgR21anKnMI1oGI4KY3rQa/4j5aVJKsYzZ6hKAnr7B96+4NJpno9WS346lYnNGPsu9/4hM
pGatiuFsYsohSLpE7l1zi4rXBtKCu/XHuElJF8g+ZTwGqMBkLn3/NKvp1aHdKpTb0J+/eu/85hBp
ZdOc5APgyYUzxiFREBlJQ1C6BYUBHaZ9PyXMxZTDQFHnduxCcl/jfLcquV/9rBZtkLfSN2odc5eK
kIeOhcHxvjVrlkRwB/2kE1yYkxdx70bIYWfEuqyRO1i2PDQ1SbNs8D/kuzb8tC8AT3J/PZd34UC2
Ku22FEtrY2kmgcFtSVX2O+LYrv1taH/hlDf+Of00zGbBF8dMU68qWQJnH1tsvRgfMXvWva0+ed3H
eSSKCzHL8PQVnf8QBy14v3MMyHD+aT+ouqZZlRfnWfvlpcAM7gr04K8kib4KA/KVquJmDiXzt7OI
mu6YGqtEik5DsFhVUNRswwzOdipnxc1Qm7ke6y3Nhyh2434J7F2o4mg/cAbwK25srPq1IanSi1jj
goRmDw3YETuXFZDruvwJTQsfgyb3Ydmx3hEaDD2zPQZBtVfzbqW37tennj9h6xsd0d+r67b91Axh
sq82SXSruF4ecysvais5JFFm19g+nvkGt7pvscWt20GQyKuqNcuLLy6RV6bvSAFC//1N6T4RrU5J
b+tmqP0XLS7Un4rxlM+8G7Ck5v4GzR7xsO5kckgZ7/KRN8IsoHZykhSnFQTRruFA1glS4jpFORqN
w2ap1xnUixa4zQHVtbbWxX20R4ye0LhBDZ4TKHhhgJ34P4ZCx6LjFiHu39TebAgYBUHCiPNnn8BK
HXGoXUycqrq6GVRbVAu84S+huFUyTmkVqO0lE9tfwIa2uZ6eDaQCnRQL4rn592sPwjdSBGyBKB3Y
BBn3P5pO0dlFm3jc/QfxnbED5Vh8FKWsPWhPMqmRhROPJ4lXCKzB4RyrK9ckfcdSygs+4Kg4nUH5
BPHFmJVq0g9WNpJSyTFdo792LLRSlbEdiLE7AX37u91Io9ljy54NTqYTxZ/ZaRAujXwOtayeyByt
HxxFUNXNG/JxHCQsiREJq5S8bRXdAGrwwhznLHZU1ALwte+xD6xKdNTGHeqg5a7Xs8SbemayaWBK
1gi3JzYiFAwT4Ui2Bb2i9mWSXiy3KN92WjhblWT90bju6jchhItnvKv0LRDKPFaJU4C27HEcQKug
JCqbX072/Ccqi0WHc9q6J3jRffXLEQCUwLBp+w1S/iuBChaGZHwL4TOLis9dap9psTngE89jKlP0
Iq3fOcRGdTmecbiIJlf2Md+SiP0zw/b2UBAukf9KHFRz0NUO+7mlAGVxt6pFerFDLWZGyLD/yERs
3cV/M0fHdMKrkmpa/C95SzEtVeIYvAw8EhPx3sg4TVHmkkx7yniAW/ETzswdreRqnsOHvZNFoLur
o6w4DLTzhEVJja1zQY4jfxp5B+zMTtQfbStYfdkPWPRtqR4fL/6slx1zPkXVYmIEhnOjWjNjDNJ3
fLfnVtMBRg1nqYjXWAnk+wFqR+fKX59MR5ZKk7NrNZnv+lqfj5nf4OPixblozvHOLVZYrjFwhGqd
siRJV3rZQSCsKcNYagB5ln+y8gVOqnN38bJGpkWLRVEyYuqK3zuIAQKztDN0U3t/8dhXlAt8RmnW
H2Iv90w6EvPuzfPijjugld9Z7bNGedDGlze+3tJbfv29YKuBbWPCPrC33Btk+nkawO0VPfAaK5z9
ZvZhqt54SFfE5I16/lhMbQ72/k1NZ48zMfrXp4ueG2Zusswv/xwGkwpJkol+sNMTKonfQfUJ9EBn
KxJ8FJSKFuRImYCqrOxpO/ackbE13/6rWHnO4QtvCpUBetyT66576jFgA+0tbjfigmUj1UxDpTp4
gG8Wthp2GaHgnfCT8zPGKgMuWMnuCJZ68gRq4bCKatDBkcuAgTb+9TT0WlJP6yK02m7xYGrowcjS
mLNeevSeZYAw90u7cmyXaqZvZIJzbpNja4GgHcCyMHK9qpFgU3nDca5qw1Da16ioTDX4KX9mm0xU
nvSjlnM6hsgBP99ket7srR0c3n/KUOijQpL+tpucLQ5K5QoVGvwrIIXag6FJqgi4oT9zYlwXqwU9
tLNJ5nxOZr4S/dsB52mTlC3egYMWv058aFuQh4KvaiX2JdjIBOoBqECXn2nNfIFtrCEwPeNhP+fH
n64Hewec+cy4TPwRy1vGSksC4kJhQXCD9wZjIxtXVOe62EZpla4qAVZq0shPekI41yPJvn+LiOBc
6cYVCjbGa8T/QX6hgzTvLzFlTY360ubZrYMQ6LcFfCmbtu+MMcwGrzg/gi0fMzcDM9wz62K4fYXH
d9TVWqQsitO9np6W4YA5glnfKwcP2ouatRLzgetbyCYmZ0Ef3Yjw32Glinv1D10qdM4iS2kIGWkX
Q/J+ydXEBdE+Wr+174IJCAmftXS+4DouJaU8dyynKFLgfsIOXh38rKHmJRNsXTiwyS5FCQJrceL9
DLN4ZXEG2LKgp06s5LKZe6kPTnYWjLoOCc5I+AVLGM73CE11u4y3nXjeEbfWksqjhqJR1Lm93Caj
9cQilEwCSCmOm7htJ2vyEnZWPpWHNeQikwQpuwdHmIoIw5oELepbAXkEcz0TOcozgd91rrwtJN0D
9jPqhCAXGSarOu3RrAlmql2eGeNnnYoFoIjW5gVrZokhjbIc5J3KF1UnutCTxOT9I123bF3iCdDd
4Ij5wNVRQnpoRuwcNjimr5o3c9wXOiSezNz4bNP2my7jSxh0RXChXmeMHnmbouOnyEBbOb9mUQ6e
2VDlG7ww0hGdym+/fEjFUjLDmX5MLmU5/p/ju0qYNda4PzDB2E2TgDKGJm94hUcARK0EoKphyLnT
CnjEYqWUxEMQM0+NNhA4zo/QH9Qm9F8Q+SL+YzOB1wVnwqupn6vyQTKGnCfPkp27MtzYkI+ztIK5
YLO8Yu4faKn2BUH24F1RW+4a7Q6XrprAmRfopVfRD3e1DnmKGfaNho9KlmZ/M2vZXrK8of+O2a0d
9NZWk4Wjl96j7SjqQdfzKQ+4Dq4oCkNzQdWUmVllY+nJ3Xy2Y7jL2KB2bi5WrNAfLYoo0E2LO+5d
Qux3f1s1V3s1bv4nH+J6Um5HibiyMcKtVEEK3yfKGKzvAq4WHpdqGm4emK+RdHnIZMd5xk04Qp87
Hr0TV1YDWLO1anbao1ddwojwlPlh/9HFcOXDIHgZULXtgwgdS+b4RllfaZ0B0iwoXmXDjfhQHDW4
YvuYMBVfc5OehqPDhG8L9QmAiArbIAMoqKDVH15jPUNVMkW3W1epwDsAeqwTErAxathnTRLM3kxw
idMzqmx59Jl4G5OiGgjq0vY31E1kNS+G48aWxkV4rFoDkRzg7lgKFcFqCEEVCf1B62X7cxB5PPSz
+bICDtW7h1AQ6vTi9vnL1or13qSLWAk03gp/HVqD++/GRDv6OimOOmQbb5uYxxRVoY2km9cxaQNk
jg8pKphHDElBnauuDCBNqZ7jvMvNIK/NP68s95DHd09c7bRtgAMaBOSU54w/Myef8kyYhr62/c7U
pxvQmF7ynXijF1Vt77ZymJlHngtbVSKe+iWaIMZ8k9DJWo5JRSsLlX3hUita3O/L9dtPABKqybyN
83N1OT7U4DyhB3r/As9fGD2dhZ7Pdi58l6oJwvUs0OFtY3n5MOtrrPElXesI9lo5/J3t+UiKry+s
EyCjCrAGE7xHh9tiLL5yfqAc2oiVw4IZTmZoZC8u4zcd4lbWvuy0JxgkpmjfIgvtL3RlivRxpPUT
kq6aUVHv4q4eUAFyGm8NA6LuygXCEumSpSv8F8pi2nrrDpvahgg/to6g5slD8SIgi5YJmHe0d5Qj
sw02hQQ+C1zP2482YBrPsT/sMRW0FcmeQiZHMob/rUhpX2wCptN2dXEED5I84v6OwlruTzZZ3RM0
G8Uhm27MEDw2u/cfPFKM0yLJy4ofOXWTRA5xi7R+m1QICOPLxuC9s9Fz1XaHf5yLqyPTEfXpyIgR
gzYKTDG35I/4Zqck0nZ3C/a3h0q5lne9Bv9htisTCt8uO8MJ87a/BTsbE7ZsibEL6e9HI8v95096
aUEggMUPxJZvfHwAvfTz0tRq7uA/QYAL5AB71eiZIEdsxYjCF7f2ozvHRebmR30BzMOSfGVanqiV
R9xG4vdkRo3WykxWp+zOACRfzG9d3EWAki3jIquNvNVCtDFPdD6nTHc7VMHeXTriDlchLoUs+yxm
tLICdCHFxLYCasrzg2fAg35Z2q9Eug0ckwzEgu/7PTbyVK4zB9RL/B5hHtCAdwAQiLOvLdwkLfhH
WVQcyCzvLXdK7bykAEP1FuMAacpb0lrQAFdJtLi4GIOrwTZ9bDiwzSjXRvDxaVmWS43hhpH+OCxO
BwKJ8WiiZVIZzHHbbZwjNVTvXbwWwDFaNxi6aj9dmg6nxIoQSecLRriE3xG7G+83sx2DttxG34as
ruCaXbSPyqDPW+oxka+epNXF7Kxg7vBRosmejfmPbaiGtLrDjQeP8bmU6qhLUU9pu4lhdG2QCybl
2nSnHXB/d42gifPwAbmOi+MELBTFoRZ5GqXWp7I6Aro8By2yeMKfiuXfrOWGiNFLMc2MJbvczxcZ
Vz5KZkpDnI3onCw9GHWNKcofb9LipQkEAjne93tGXPLIlBzn0dZSP1+u8hXiuD+VFEHsi3KZIMZi
f+FBg4nSW6mrUSHewdbaQS723YVWm3HW7NlT3E2dQFDiEiDsEYoL+lbmFTW7ko70jyFZ/up1kYM9
KzxN8mFPMZjqT32sMojH9A2L+d/KBTOGA1fJm2LLnPCyydOLGWjLDD5iyRn4jEI5IvWInkbWOGGD
DoWmPabxYK3UWJuLjUO51YmQKYAAPJDeliCkykBH5VVtcO2KwjoskrqxdrmZ1S2JzTAMmCnCiD1W
JIfVnv4TJgDIrillSAlFCqEDx8RiMc0hkktAYwA38R2evhf0Dh0iOAdoaJuybb1P8BCWF+MReMwI
gCXlX0LsewMQ3aBqTwVGlxWhfbxy1R7uz1sSA/mfE+lvT0FAjegQzEiP3xaUz2ZNAbl7g3zLOUi7
2VVKa4uPo+um1UVNgNv6In2T/0wo6HPuaRmqCLfe1ibraZVc1VCRN5Qy2mXOGkKRgW105UyfATOm
V0tvvROskYMM/23XDsn4DrJNTwfw1CwFZVAtRdDPsnpPSVGI5C42Gz2L511/GVU6Sq5tMNjZQ9JJ
1a8+m9othaOKzBd0FY8SJtLbrN5FjhlUOEhSw1cFVUaUwFT8P6XG6SXeG92moKb9GIUCZ/5Gve04
1tAoiCq+Nc4/PX6Oe81XahmtLCfHo5txAY2hzvZ2/QIdDxdq1oOe1I5OB10BaT6SOb6+i7yW7l0S
s/tGKtvkkMk9OHfo1NW95TStIA6f1jg43fZvEx3Bx2yyeAoTF1pNIKa4EXXs8USW9c0iG4k/EmDq
tLIrEsWB/NQuv13VPFkBeVq0weloED6EbJ/XhDThLxvvWCFeEqz5JHLGHPq6M4FLIhPfUGlLEsGC
Kwtv8Uin3uUecnJKi0HlyTQaKFt4XK4205aZ4CAz3ON2E+gxwi6lqL3a76kaUsSXBD2O4GuEDNv0
WhDSKacXpj6DxAxgxk57+cQNjNQ/g/wJVpTN2KQQM3E2X5nC2IDWDtbWYCfTylGrinps6pOEvryg
dMVJNFjgbs6ZtUsOXcirZn3P1UMe1srsr12jSRPg5xQfC240lW9mGknu3TDz38D4XvdHLAVpcqNR
u8CwKrin8ZB43z1D88B7THI0Be6S87EIJGFNZarMn1R8oUeiwZAXIhXSGV51psjXjXiEZ4gfSWR2
2Ng6YXZOmkDWIOijVbEzEE5w0RTkvFQrh3LcopThvvFGTwx0DgkmQbjigvBpOhZ7iwnOezVjIrMP
O9hI42pdtZVoiagTNTVyeczgAdrcevcOQVYoOylgHu2/MSL1+kEafhiUIxTYah8tNNcUNRbNHjas
OPyScDikmQW+rFbzgNU+mrQHUoDyFDplIAOFr4utW2KwaHk4+5QoERoGJZ94Bau10yrlslIQxrSR
1//ObFQhzgF23YaXhXyg+rCnbiXhfb+WH4GL1jBLZdvK7lWrFEUjDm1j712d4FaSMTp9WC47FuKm
VgrjkrjS7vTJnbirTSnK6+Cb/5gt6udDAGego0re4DzFiks19E42B7z0WMCJbOJcnxrDXApv/8JS
VSeH1hZEzTi3Cnwe6pkyC60fOZM/XzNqNfhyJsP8sRR5E4DEBQgMTYI6NHudn7MfStKqaMProN1b
8HhbvkEwjJgLHMMp7V50sQkuMH8fetmiJio8rCM0slQ+YZ/U9dOW9TT3uUPAPrKGoB2q+ez/o7lh
LsEuaeALk/Pit8X247RNY99gcEzUjXmtzKeoBtNpn1fBYk3r6qETneTIDnVT3HqjwnnVxFi5gLiV
IUOXqvdDJt6/DKr60AzlVQwD9ChvHvJuUwZ70U5buepxpJ+/8MmQ7UXyE/5lON5/EGxv1qE66ebe
ZLZXcr5rWGv8PcKZgnSlq8c4wLgeMQE0gf+etV2naB89uYduJI01QBpQtpcoapfCHjWJiELlnooz
6BmlYTx7pyI/3TBj88jwQUfvWSDdxUdBmApj8/AhSw5wpnFDLApOoSM4QjOYXczOD5mjewZTaqEm
rbkNDM6mCAkbMhg7WXsKlgLQi4kz4XoZuYj+gqI7mgTFcc/HdhZDyCGX+oeJX2CGXDYAQjEs6QNe
JdTMnULQ8iPrWTo8oc+E2fs3Uj0i4K392OEzx2qjrkdKDtyHCuWhIkrndZl+uqqzkPQr3HfW8Nck
VhOLze8dH8/B0VdOyMGRITGh+JimmWs4Jg/JA1E8PdPeSF1BEk+H8b/rYHkN1YLz3kJtR38RzQah
ilgz/Q4HQjpo3i4dUxmBASllyRhxq1djpwX9rtm9+UqJYq5rJB0RwFS7IhrKwEZNqkhiSFciODJM
BEJiKRMkJBllXfUXAcW9HT5tO4zeCE+rZ+1NYmIfupb7A3q8Su8pEHlhG5HrUMvK5oy0yLKyLqLM
KBLnTbgAsFoGnn1MLvePt0jcLQhrCuIrvdA9sYBjiKlPesU9s0CBjVSj3YvYzB5I10zw0xxVqNZC
dIaWztiRQ3A6yCoGIOq0TKfZgiKKF2d5oXhFucO+JKfiZRY4V1M4Uzt1IQR8+4154rADMlNCnI+j
uOZRSfsbvrCtEKyuhnv+PU7BvMPInmZz0Ing/MgzFrvNKL5KvsAnoNrQTOoX+CSbYEyQYRIkdOPO
67bXY6ghBIxBgkuwUP3QV+n3r8VCCCC9WPwKpKOKE6B4Ovu6hTgtPDIzwyEs9K3jLHwCpaJ5/TcV
atEVDEwilZkmIKOK4vvkChkYTjVlzfUu4aeSHGyeZXRHZRlcJY5U5u7JUZiZtfc0KPKZLzXfh9RO
8gfA0bqlg55ca5eBy1VYS+wLJi2k3tX/Dw8vLST8qFdni/4IXNFEo+rKgmfWPvY9/cHRZW5PCeAm
b2fv9nlIV4MBEekUPdWNoeUQEEHJiO+ODo3C13xhbqytfcbCrdJoHl9W2zApQ2Lorc4yq3HIIlKS
vIRoV/T+A8SIqXexI6BbYm48bzj/Evu58TrINTB1Bv2LvVxRw+Mf18RUtwjYIlp01fU9zR0mqki8
etXjQ+SMAvD98HuI1NdM4CdrlMcPxh/jQoztluU8jFFDfzpVENoRQvSZGykvD8MKN7Gjq31XTh7s
RJOXN1ZRFDDKf0QCXr9sKaPgvwZMJDDW38EPmRcEasT14hcpGbjcecs/f01qVpYFJQj2V4uJbd61
ChsjZj6EP3JJuEP6Z0xAT1x4DP8UrXy/eQIBtrE9R07FE4zh+xbEILDj0oMSRNbbwFnMBwBIGFWK
2+ljOwziAEs2LJUaUfEhvizIEbR491VtGG1xbt/1IsBU8stxAVKfxpTJE0MC0qMkmkZ/d39br8iu
BlZrhSck3pbPpk/c249WxwkmslaufNmqbDUXjRahY6i5ycoE6KJ3exLizZYfingX83Xih7BH12vr
vF1iOfAkqApCah03qU9zrhtPnyFBxx/hao09+WrmhE3xPw+QSslw2Zl5fos6JwLKraxDF9swWq8N
cEGRQ87Ps4NWfHEAzRTYRE5fM+ZfEup4pW44tkvk/bHJoXNhSGxOIgdl3pwWQOp6HjSWdernQyPt
cXIpZ5PiRyVJIU1Q61pUmG45T8Jxd7w5eJxQwx7WFvTKZdnXepa2HbgYf+pPo875UzDaQCFNcuKp
UIHjpSvsACzGO9UA8p2UnT0wuYWApB1vyaiv4qGrrZsC9LPutdZQTPxorG6DXundvpWyjqbbj2Uy
moKrpiKBOzwg9UHc+zw7PIdheT+GUFCA3ehqOJ7T41LkNdjlD4t1Enl+0OV3mZnNjKGRmRlArhCT
wBsUkRt7Qvlu/FJr3oJY/6yOo0bJcBwY6h0+Xx03UxgXiLDuO/h5foIN2A94u0dlBmfNC94+4Rd/
2IwahFuj53FiTkr9teVAcnw1U+UUOmLwtZo7KJdIiEM+c6QKTYzEk9Z47S9voGwZuymwXkfWgWsy
ffRp0lo4LWBYZETc29oe7kmq1BREodDpJiCyTUSiY9pEFoX2Q1fefItZmVIC/C6N8KfLDcun1Zy4
ThWNk0KkpfSuvuDvyCRBGMfOI/IvcLaE4Olf/vEI/FKsKj72kNQrlsCP951E6dbJyt7o2/9SMxb1
/nXUJvEruJsC844GX04TtuhZja0LIVBBcgr2Yde0nk5lBrDkJpsG7C92As6s2/6bbH+IV7CCaxjH
EPMoqslooZiYyZYVgGOePPUYniMiMeV//wW/Zyfqmee2/lscTWo0fa66U4Kol/Ih4MMoWfnYDnGC
5ESg8WQAxlGpQsEQxzkC1Ar9sxfYIaF4N16xTfZ65t6PX2h62hOTTueHnEsDCy17vfm5TMUZOeHn
aNXteKWAOM2g4AATgekMS3IEco4Q+Y/YvvRybcO6IlCh5habs+bIe6phl3QhF2h1EtfJY2gUTwfM
CpBEhwOsOn78OvruiO3eP/qv18n13RfEcvB7dB9qhcpPMupqnWbut5pFzCr+Y/5elKR09dtxjkmD
DdDD0rBe2iRBSUn5QlqkpIhJKmkViOKw9hDZrRfdFOvxW3/qzL+3O7/1a+g6LJYrsjARVirZBIpt
bJ4bZTMp7HQsRVqaIQIsdt36ZK6427N1cKwPfxKG42SELOrWIjtvt1DtZ5X6C3JduxL8ORxzmb9M
6tOVm8/s86qvghv+Pnqta3/7LXUiju4VsaHZ8cSXmBDi5++bhT5e5z65W/sHJ4Xb19zTNFaf9Cq/
uxAnMC3hD73p9Y2hWsxdrA+CyNTD/MtrMw0M5535QwprdjAvpiTGY+0oElPzZhz11f0s7MPJIhTP
kSNXcF1B4jkmaxeiBJUoZyGdBU9Kz+U+thaQorMfyvsgEYeTtd6vho03olxDktAbU7MTYO+WcIzC
h6Tq3FCi5U4H2CVY2SX2Uz6O2lkjV7K/xPKQYbARiezgmkS7BOOrgZkwEywvMjz774yVnqRge4xH
8VNHXTUifH8MINClgDW+nvLMt3GKvFsPNGj4FY8MSmqb3rZ8uxkRVCoWs92aD0xwnnJhQHNSkhYE
dLj5bkRakkee831vFzRhETLNRktYBaA+E+20y5ZYYbmiSSDU/dtLYQDwVI8n00w7bDaw3Q1AThLZ
I/6VQVH1qlhgnqb48KNJAV7+hJaQhG8zY0KyJG+HUrjhRLb77BANgIOgD9JAnMY/g3hkiLDrLtwo
1MF0mW7MRgjByoHj3juFh5IeFVzliQNQxWrOHh080J70aVq/knqJlqskcVyoenkU2oTntRDAgq2n
heYZvKkeiS8b0k/04/Y+HYu7+Dd9TN6sis2xMIKyIMM3cOIa57SvSP0d1aSqgypufWE6yagOeViV
gb/FJcwtTtfOIXoeaXX0i2aUNSP8EYwLFeakuMnVmomGpjCzdhCeuC/aZmpNtVLZ1hX1S/HvJ1Zs
SOmHuX09ifGTx03XBhdML08k570HbkOnTP+cmzzslqYz2PtDJ5jEKYm0mrz7Nhzy96Y2KaH0/syw
IvZkJejebeFXAkgE+Xn4/Zr7pL53Is0Zmrk2hq/TsiDoDLT9/ZgYbyNWue9Tc7gaD4FwV2cLAFec
NnfMveu3KikWyu+M3CclsoFWJTMrnBieCyCWK3o6cu8yNQg0nmZUDsjBq94McmwWPvMLj1Ezm7Lw
cexLmuqLXOW4RWj+UVI4LooPR3dc0rh37dbXf5irwL+IiUFaK93b6c0lA8tmoWQFf9Cf00508AN8
5J9ovr3E0fzX8hUCZoIFYMlhQJnIcmr0/7kEfTjMiCRHo+pg8mHrqRj4aWb19Gbe5Ngx3ZQZK74l
qdbDv3n7p3vB8M7b3uzUVK5zVZR3P8wdpP6km9d381TQvVdaRrFPjQJe1ew62c24b3RuRPk5BoXH
IEXJCeHzA8CXpZKmM2EUXPGn4vJWO9hcIIBKra2PHayBnOIG+P08vhQBafERkvfWLIZdOHM1KX93
iAomwSYGZNb1E+CjKKyGfJPeBLw8s9OmSde4Fb+CZ41rtMWDWssunjEjbtFOsWZ63g0xy2yZo35+
+VTGzO+6h73V5IFCsRdFM+ppqyjExsr/aDrR2lwvWDlmHwH5OrPiHv418OzrMT2i2RU98ENWbToY
8uH2lJ5WXfhjIR3yqAuGOOairbSTl9YiQ0BPSD3qXJTdqNwV4hjKLAdnyFRC4WkUgzjFdNhcHxdY
JC9/FNE8v0EUZM3hO+BR0tAl5io3Ld1PCszinLz8r4XbtxTrd/Ej8AZI8wg0GZF6PPmWbQ3hihsR
me/g1WcQ8i32kFfK2CmITYbOgOEQngp7L06NWAdqD8JlI7rFpctMeB0yxq1YHA7Gb7+nNsMbezMz
zWCPfLYaFaSc5DUOSHIno4jjJBiPyKiD++EJJUkrHhL/CgCeOstWyXWSTbkA9HJgV68FZzP8jvxh
ewl3fGt66TK9OZpDt+dg3ymlXoa50mPz1Ds8Wsuzv8/eD0igFRHG10ItYYt0I+dbZZa9jcglvXWr
LXMbO9zEXYLuClshbiGl8Ae8AdIgynKcXXbjVKGR1aeM9o12QuTfP8ufD4C2WBGJMLNfSuPzONy5
6EmRkbxFdpsM1xWfRZhOYmEs/UhfqY/RRuuwlw+u2K8Md6Uof/NWjIe/MUUB/nzgiBboObw1cIED
54+cc32yII6XKXCW7R0vXjnwL5xu2nfX3JD63Ul0Eo8dRUlQqvmAdkShW91TCZBIqW44BnQzUwQk
B0sw5kv4Fez2AHQL1kijoR3LEhAN6G+8w7JBt9LyKJ58djRrriELOA8WSA02XveZvsiBtAL60HMp
AICAmjWBN1oqL3f6JD+KiaHlvmLyWOx0pR37yqHysQXClmjYldaJ/HaOT8xBEKYCvGCKbyBowSPV
HzBenotUYnFYgzuS7rsIaceYro8apnTU12jQsDV2KNMcNrijbk/+BFcZJjYvPVkEkqFuTT02s4Lu
NKCVSKU1onDQ+i0Lm9gdkEGoMlEKsu19mxme82Yz/WmF1GS46fONVJPcOQNAO+DNNEVn0ZBjbzLb
P+IFAeKLoZEHqvLBsRyube149GGmBe57hID9qRtiM0Te5V+kBccTm0i509TSnY3PsqJaTEcBgBZv
G8T6N4b7G/dcRte/hKweq7pWqZFzyEFKGPHH/7uZ9VlMiXf6wvqoh0KcThCj/1+XMEpZcKfS0FFB
w6s00AtihZ8dCoJA8KZN8pZGjE07kqT85u0kmlFnuFLpiqUH8CTxzeVRStVI7Xhq99qrkZ/d2xtX
qdXyKPYBNuKsEERwYXZYyfvhfSB/+w2/VMN6RmkvEVr+71USiARmskpJYEhajc5xkkNe+4Jcbc5u
c2Rg8gMnmuBvA4Ad7zJ2NgvKqi8sEgRnWovOr3TVh61tDh5MxvgX1cXp/5CetsxB1DJYocufxU5w
GZZQrFUrEqm+oWcY4MZJE/7vTIO7iTTtG+mMsMnNYhWH49KqM6neIX2R4CtMm/jELnIhoF6+t5Bv
OS46bRIQtv90naUKebmU3R/hRFmC4YrApHwgiB1LsUjSS60F26vsUAxMhBbBI71H/NYK2Wlntu21
bP18a4Q8alm+H6Kwq4ficmLjrIx6vbXiWLX61ClXS/VerAmMjFCt6P0G0Cz+S9IX/nrg57WMlH+S
DTamct+HcDauRSSRJucpPq5rUinWL/MNKudeyObDbTh47dyttR7Fau38A9SgjOe+rZWw345J0IA+
kNJyHGHWwcxIOBa+q+QYHvqfDvYdc69QffPf+5Px3+zy2GN7QkedE5kuW8yyTSd1ABAHL5ecXKHo
4LJPVfc1w9/zCPO5tnlF8wvUIZzTD/p+wjLAmVJQcnOJVyluCsUp6up2Sz6UVNu+YvENfxV1angW
h7UnLY96J0mVeXbzJbVM4WtTZ9zeuCk8glasbOnD/FCH5p5cZ7kU4oZjUkroCIvZNboghGvvw8XJ
3kU+Lkox1Kc2+B7vQBH+QOZUdhbWYMQowSHDOoaH3DudqNhanvKpHsWm7+GbCyj4jDavB6rD0YzQ
XepDu9BmJiKNlJmaLWu7Jw76yALO546lQ9/xb0/ox/IN9mXpCo823ZvfqojGSWrTv0JaI2veqCSY
ZxyrpvuXIDD6wYvpQ1btX9hZYkPepZgSMB7kilauYHDcXPIxMuSTmf/M/5M/CWxoW9V3o07CNqNp
LlLMVuy1bVv1Dgg2oecczuxzbZuUsB1VQ4cBFXjiDll2phpj65btCPsBtZrIcxIBO/IIw8ZUifGe
guCFno7IXlFp5y+O1tTK7No5PnsrGYgRisNhFWck/0PdoZEIZ9VR9FywaI0M9taw1/wmsQgHx3tl
cxSb5PFeCv3UgTr7x6K5yR9jGH6Fn7DUHhOrKCX+zsTd1hdmJktbdzOGVD9YE28pOYqx+4l7dZ6v
TxHzUgCgwrb8wGOmcNT70npxQEQQ8jAwzkS21FAmZYfxqpm+QxPjeWgiF3feRXxFCKXhnFRcpkbp
4D1KsrmGU0fccWqHI0j5h0PIPeeoJiHWubxaEWxHF0blWDSMgOqPndGI+cos5aLPCShqj4/fQCO+
hP+nSJ0X6Zwa/Us0o64YaVHrdv/QOnYOlZtIXQbmr0WRvmjmdAcqd/WyapV8bOcEq+i025NxF0zI
PuRZI4R3aXZyOqz2TH3W2uCeb7SVyhTWHs/CHSIdvf/jpA9L8csS3he4JvFlfY3wWDTQA7JuOURN
9Roj5EE1IUFtNY5DB6X5DKC4l5V2H1XB2j43BMZ+1eXH9GWKHJAFG/D5mmtSD+d7cpk2BIx38QX9
y4qjlnqbqVEG89VEr0c/L4DzN+kP5N3TGt37e3zba4iGxs1rbDwbylCrFDER94iCrAfGxGFcfVOX
icd+J8jj0AxxDYOHfa0wGSOp5G3pi7/M3+My4ZY/aV5Q/KOHUQMOI//JNbGSKcPGDVVgtffZg1zK
2nTGUEFUcPjJRrw0Rlq6sND3touIg0j2NKfaJwG9g5QO40FzgicNY3EdZftQxn/ZHj86Vm4fBnv9
XYknuC+ylKwflDiQYdKnYrmH6pcoVWZZIpC29MgLMk1eYTCm5wf00sevpY6BVScLy/Z4rAt8sWEc
H36uw1RdiseHXmV379ujcEpsmHoSC56kMLgaro7xqcwHFJo7Z4TUb6zyiiGxF8H9NC08ngk72quj
rOQ8dXobC9hHnMnJSzHuHTTgQNlHDcqbExWnABX6lAapVbIuHpRjoOPIUHKeQ5B4adjRy8ZeF6FX
z/5xsNQ/RGA6Ynp6bT5tCMKnJ0WzULvfDMkz6C1n/ZNl6HHmP3eIF89j0SuvpGjiDqaBY3jgYKQj
KChrf2kfnvDsiCwLWGjW97BVVVg533hiMgACzOrF9139Dh8k4EFPA6eLlUM9KwHd8rExmSNU3coY
bajdyyawJPo7D/Sq4wzdTxKV1FQWo2hJk3Jq1OoU1sNLPVm5XizbUD2t64q7YEC5wFSkKnAr51xX
eaHZXqup9+et3rRYLVBa6vIGeWiPDorfpZoKCW+Q3oEPoHHdINJOxarwRBRf+jnjL4A/WRvNcpYZ
V5NX1sEoTpNf5LcNLccKsCNBkedCXfMcbgR1O93BR/xp/DBHpOyJTiDsXWAZXH4oW0Ui8Pb6hvqp
xlP7YO+XHFXXyzOIEeYZYxY/1ceQI0Vdp81jySXE98kx2xUQ1LGQZ3tSuK52q+TZc1sYb8m0wN0G
U0ukbnlkychOIF+ZCXuZSXeaxQ/yQFrfdYi3m46vKpbsSBi/MxZA3CUpJ6sc4bUPtWmS90iqW4U6
B7Ys3FyTG8XrBaBYJkg+GiqVlmOrrGZC49iMbhrh4KkjGtOEI6D/09pYOqB5kweIgddxDbElYUH4
X+94ptgIM3QIl3jkbwAynwCNXy0OAVxsJgOe0lCDXTuC7qcO6aSvGScptfgpoXCoN4beBHuLOIzC
tbbfWsXlst5tkPPaYgxoetoc807mPgrVoKyWkCDYQgaFTaDINvdlZJ76NLwWLMbzflhGMVWei1uS
pZml16ezGZwKVK8lVJSOPoRWAwvnJ8rBcnqy3w5HMBN59QQzXJNiS/S2v0xTafh39glSfypBSJMP
kvi84yBFP3hH8XvI2XvuYYENTQE15R6W9GIAz/ChBy1C9sBxkSF7xh0BWS7jmpmsJ7KkrBb21R/a
GF1xC0tmAyrKe/qbMQPnMN/IGu3RwYrEX+B/vsyxazqkqYWlrsCu74CUVpiDBkV1bEO0/84ulRBt
a1KK6UrHzby6CspLpC2r1cVbpFsVOhTSj/Q4RxkFxl+HtTqkxA+lbIy9i7bz1yO30E+0MHAlI5yp
ClS+GzYPukXWkoc54B2H6vlVIPQCXXxkxrorAGSo3rJnaT/WMzSjko1pmMONWF1tywaIXfTTYPXD
lEj8NEfRSKbE/yFW6glu0qFBhakKByJ59I+TdLLxgNKXkCDd84XLTC5nm36GCVPywxY5PYT4f0EB
kn4oQo5X+MOczeihlozBx3OVX+vhyyeMvSb5R60WOIsupY6LcnRstRWgPjwETCShffcdEKvFJYRp
eCp7Mk3GUM8AVhwbPsF5dHfjf3JmAKZSdlWR0K7GCXnH/kVSXNReAB2Ff3rGQX7VQryPOW2TgURU
uQ136l8Q/nYQuEKnhedePOQBOH34ladxYb8b5cgjw/e4EKetc5rLyyittFOPwSKapq7WGzP0TamR
EVaV0ypjCZJvwwk/ESdx0Kq4IKjklD3V1pq4Z7KDqTYBraa61UK4Fsvilghd9Jy8VCo1j8TGem6F
jydFhPFmnkYB+s5szfAxu3PcfFKH4T0/EMN27TPJlxxFL/TmHdCHnFklhLdWc075vdKzR/GsgPR7
7nSjfwJrlUh44eIHEzA9LqgpEUavtkb+vCIji6b+a/t3AFL7kBO+gxrbkHYKUoQLAMFJbUmyLX5U
naVnoqMDC6s0yGZjKYBIb7N6BedvUqLiodH2gRQa5T7p3wj/vqltz/w5NuM4Iq1k8Kr3R6AyydlU
w1S4EP9GI5jHl2IRnKMJgEV/JdLoyY52ZhZ4dfnoeXgO+Hq0Y2YkaOXYhtw6LmJZWmFA+OwlfWzJ
ZBhfiWnRaUtaK+vhqouaN6qwzlgWjgk4xndiShiiZ5KwbTFNjn2PUoVAcTh8AR1Q04/UBy35Grdk
icOkq0CMYeuF7zBz73CxPDZSIQ03rES6cETVYwuwariMUot9SAiYPB+NzWCC/z+gZPKkjxOR3lzW
I1WBbahx547g3Vm63rQHB8g08xp8xfjIS3QKFEA+GObeKCr4Iz2bPVa5XY00cYj2JndA3idurlzk
It+SuZyMQwHfPGV9P8B9WTQ0qpnEybq2RBi/uuClO7lRi/nskWeNHkdDOAHim8oSl+LCVizcaaK7
Xil5PpwfT9rbtoEWKvY1C1hfCVda/inzlAGGTDL+Jd8PqzhX0Sn+Io5sbA377xd8WjAipxhoPyuT
az05DViaq5L5BaBXi6QZEXNI0hJ7xuMzg2gwnyJpgmp+SK8nR3PFgYPz7ZcGANq9/0wCyrp/LXrw
zbwCuxrBE3P1QGcsZ4uSKQmRRrvKB4lOqGOmPHKzC8lNrHxuGgMyKIjIrszLfMBGJKQBULZqcrVm
FsayMDCyw1woTmo03dYKw1a3McxD3gJFTQItaGKxV+FqaGsxVmRVycuU3Xha45u3tfoCdaOYQzrI
UZ/XzeuoEfDCxGW+4u8x2Z9K+BZQTG87TX5rEO/b9ei1Das/zSB+b40SlAB1UzsrRaeVeL+GyHR7
qauIS6JDe7dpU4LCYevBcZBFz5iMuJFOM9njSsn02+4W3d+n/aaKmRP6YU6hjsl04+Hjzo2sVFgQ
39TGKHzN2VnCLWTVnujn0vOxU+vKumnAt8e0B1o+78TUv/5H0f9t66Kdf8h/u9Pqv02oyfU1qI/I
/pFU+2w7ErtpwYTuGvC6/Ba+qEmZ24/Ktx2ytIOk7nTS8w8e1zx183EY0uFI7IMrsyBaMt4NGJJE
28HIDSL+yrCqm4KbJ9toOpwvMs5rwf1rmv6Zl4x2oriF9lb9xqa+Wiv4Dfs/nC4KIE+Z4AAiKoRf
lGJM3JORKu4E7rk3qq3vKpqSARv/Cehb4mSAvTvbkh4Kzinxa6ub/Gpehw8VaPhsOtxTMv07q5oE
0g9KT7s0XIEf4aQxxruqnp7M4AzIVVNkPAHJH3ggAIaYS8iGKYt9splDvNE4mTSENt/OXY5KSoEM
fE5Qku0eCVcWS7nbUJouhtY7HKtg3PzRPGRFak+WTX31MAV7freHD9f+mne1GMxUegrGIpAwzzC8
uN3TpLMtUlyq78LviQym6NQMIYq1Byo8ToXDaru/FBao/isKOil5+JT+/qECk07PBY87yu3Kvsji
ky9wmhkyfobZ7dOnPEQEyo31z8Np3su1Ex3c8EdFqmYR0J6hfUZKwKOZQweLFJzqxZb5bpCP7b06
T3jniDVowhpVfseggwrt2bNGOa/a0Id5LlI4FE42Qduj/ay4Vo6cNtoVMDDuQ3Xk5xKlY426/ROj
BP9Qpai3h61RbmhKLOLqiIjPGrHQUkw2MjNPMbkhz25yLl0liqJAJIvLIXiY3NOfUbrFNorzkPD7
MiMF0ukPWS9ada0RNC7xb+l3eR0Oqn+ekYuadip1OoFJ6DKOH8NlhzezSYo5rEo/78sXMUwo4una
t1LQLWdrdd5a7cjZbCw0dX84qt0RRfbNC+OnRwGuM/pPTZMhGDR6bTz1QQlvuXO1qs8TGs/Xk0km
2e/Vl+G3PQLL8JGSDY2p6hEna6rq0bAX4ciQNz5PLqzNO8PWL7638s4pXRQzOgBHyXU2Ux6yOOH4
x+4xtF/MJNKfHSKJBg0xmy5aWkdVg/mAa3KDnvB2oFfXXiWSwvQMrAl8HgXWG9D8VZAJWzJFFdKU
UxtLPR4em9Qyv4ts1wmbXJpQgds9dAoPpfi9lwMz45ithu6F/sqBY49+4VWgNhB3H0ahs5sUhLmg
gwcklNjh4FP0JlZk6wJvERBe+5CNAL5gRv3zPi5IWoo2rbY34J4JWCzgQdOTJ9AcEBJEq3oI6fnr
aknvB/eL/xeQLJEXwNlcHQZNiPV+QxSgevKvjpxJtfFcdjS7aTJjQTSB0tt/8T4PDiiu1+EQ17ox
L616FEqmeoXQGUFHHud/M7Eq/VFWLJnvtzq0T7RL2+PV0fclzOTcDO3EpwugF7GIbq10nErzzNwp
vtNbJe/xRxs6UG0xkbz2oRA02p6Q0yHvMn5gNJsneYak5oEKp4k/W/pbArIpBvpcqbZCuvlaVnBq
EO6Au26yiagmPW4SFt4uWC6WPoidnEsYFaVAue4V5k+742japrA7PNR08IdbwnWOntUOydDOJa4u
vBEJ6MGaC6orcA0boWpKg+/r1WE6XrwkYacEXJMkpzgt2U4oXTvZjr8G6lYfv1p+pCYVAX0BMrbA
M0FQc5+4zuXfkwk4hiq07WRMDkV09nD34j78IBXUWMLRf8HEzcEKfg5nxbfGWd3omqAVzpeFkLDP
+PEHGAx5BBfspyGE9Q54shH0o0e8GqshDv3OE+RWAvv+dpymlr7M7iVeDKiWK5eXOztoNLA73ntV
+gNnZfR5kq/c8qifHLuwd+yKIdXJEhiIYwRCxiU90UiTalqevUTre7/kM5OVzgAK6xA0Izzg1g6l
t/FL0hGnn0AU4XrBjFgjcJxMKfxBR4dV1Ptpm+zzrYSqG/HAYXekwnvEcpKYhAQaJqcuKYrRbiFe
HLMCnV/D6QQKG//cwdMgmKQZ+KR451Lt5BJBX+m8KmIrFGo1uVymCm45W+yxcDt0igOa92EgclSn
oZiiVOyVZvRX/6txJU1+wntXntNWj2g59UyYpEI4mJBTj4EMIUp/H4gU8YRQOJ8JAX0R7b+H6l8r
AuXbsyFAEG68emMbvMh3RU6UIMWSmrcN6euYNCvxFfoE/ChSpiPg5NuQ35+Fjb2E6PUKf8854xKV
MIrNuw9Uex7owRV5Xv3QO6vW7CsM0moPTZOIz/yp60JPoPYFbYnu+u+vGY1fM5JfHSgbOQQp2owl
NQZkOW8iITCNqyAexB4qerSQpF8vyxmRnXRfOfddkn29vkEj9ARyzLlykA5DSiQtJKq7fYMX4pVl
mr/+mEpkFxKI9HbiwB12tDjWL9AHqKiwzTa8KV1sFRCm+mlQmY11CHckrmWAbAQMuFTok4dqtbf6
ng4G9MdWKytbhEomKv17ab6Kw2VVBgbUZONUfuycQA3ZQIPHH5qmVdV4RdMwhIluFKM/sFc/onZL
mHf70ANJr3FKpC4x/35Mmm51UDTP6sZsTwLaw6cKgr6hNwQ2YgEEVxP19lCtM9DVrl9CQ2hLxnKN
3vhRt9QT3tl+KRr0P/5axdrPfuhPHlEIif+HBbH5zYV9t+3PilyeJliUupsYzYN+5q6uQu4iYgMT
eS4lEynCUJEe1xfdCHuDsH1kiB6Bs7BZ1gC+D8yyUhUqZn4IJ3OO8VH9rK8VSQmAhUVRmGmZXTu1
3PTpQsFIugf1FJmB+iMbi5r9M8DX7jd33s/iaPWQWyo6gAPWqoxmJTEgiN7XlEDc83aKNG5+pDOU
tTbXkR80skKo9wK7sZlWQvfyDxrTvGYqnuNv1e5lJ0SChkskpe6oZVnxWw0kGih9DJOCpd6pNFX6
HTQop4PZI2Yko2wV9HEQI73YKHteuvP5UcUpII00XOxZeegUe+H2WdtKnUIFGd3WEdzPUtwQf6p2
5OeYA3NXiA8n2oiAlkoHc6T+im/Fudcx7HdNcQ0jqlNV1TZUML/Oz2WIwRh3bgEOEcfIWDELIbEO
gGk77Py5Z4rr0NNsoFurgD2spUCO6y6fd3j4GuGcEtG9AzKRK17bMFYzzW+ibPcQ6HgMrx7VhIGH
cYxturCnuMr+caE7fZbBVmvvfO348KchhvrdP9SJAvXS2QIuXJOUTqaxjkv1ApEitTk4zVLJdHzf
sVjXaNOELkHVS6LXWR+F6I1m21oZ16tcAX1iADEnDCv2heOaSH07dL0EdTOfWXvm9vGoR4i5XXCD
WaANLCKJzenOYxntWQz1QZZQiYeMhnNmKowuiQKbsTJbgURUQ8/QQogifYbfkkMk7sqmP8vchBQv
05Cx8A/JKTWaxL+pGknKP6AohZZiKYp/SykQo5KuyTmNkaX6t6pEj9m/P7zXeeb+B4Ir6WuH0KGJ
W4Zi2fh6vhsw5MoPe1751z7Z8xyI1Egtqcd4XAWLtSfOtpzGUFpiHhXAwb+CpIc7wr68SCiAW58e
vkWA+NSTi4Q7UOADO1CQxUhvG784fHQ8nXTi4OVBwJzAQ0w274kEOsdIb8hGBDdXTvLxJXvLRD5E
4kW/k7Lx9mNeI1NAYWenWfmrW615BDW1tsh+F0JhLuEGphbbbXb2zGn64zrHDaDC6Hdp3onhl5Jn
WQYH02Bv+d2sR1JLrVIG3VT9PAb63rJheshdWwXngndECE9lLbzTiiNvkrYDOI7In1aEV74H+J4l
a3ZVIG/zcRHROdbwNxo/e/2NJk5HhtF8Vw4lBneLTEUZEUzZEno7gsR3KeBsdN5MHPOymCUeKlRv
9HG8CMaAxxfNW19YVOGqVviaCZeZrjAIBpg+4WKqXiVLdwc/Y1T3sPxXG42+XFXJAyBtdU4j+Vz5
/fh4Ha0f3IS74Dwv2Vivt04rZB5g9ParqDjO+0U9EOVWGrwrsvMBByWaj4KXK3hfkCF/M0nyaCsH
3pnGZBF9VacapOVUHxzm9pH+UNI83++422zoQR/U9irCgKizpEVt0aeYPsl/lCumgkYzH9z7QHK4
4Diz3gRGJzKH6aoJABfyGs9jfY7dNtHu8UZ3K503DKOyJOnBRoMwDC88WeLBQ5/W7RodNGQZ5vob
uMhOHoVPdgcw2wj+cx+yB0n0svkrKJm2zLm1r+J/RRBTIfUN8rCewJ7Um01Zo6Yr8h0jLxJ4CnXb
zqCq6BpWTIX3LMqUBUdsHU2pzVBcfo/VnmbdCan8Iw17ReK01mcyuuNW8nU+Vece7qyR3y6ghsWt
wYbVvI3e9kO1rzuVH89pPAzwt1NIUcqXTyGreyIvHeTG6gluLgrKnW402Eqop4UDwq0HfHby0ijf
JFl2/UUz75NLQGUH0k0D+vtSNaw1q6l8PX/D1KQLZwF82tZZd9zwiDekrzMo9hAWwSeyR7Nzz/Qx
VpDEFwNK2Umeg+DGh9iTzLCgreiMyiNlwNdI+cc+SLO9cyzhSehfnWbb6Q1pUw9bWF0Lp4/zpYN8
fhOJo5SLqhq9hd2SkwjQrLPZIeWWdRiG3b6qZeAHkztvOUZe/2JzoQEj6jSayGnnFSUj23I+rqME
CP9D9j/Ly4dEckTqB4nMEzaSeFAJKOzOaBBqs3sjUtlZyPb7NKRZirMKG/d/iKwE3norlU9NSjFo
4gcoBB9ciEaTiDzQ7DPaGCOxAi8wSaShMo05ULPcYgcuy8p86OgeiOi+JjrNSAP+s+DlhpUm++sQ
O/W6RhUhjFqC0xzYaF83VXr5LUW8mEMiewpMJrTbfO+cyn1Mxfn7IalnObPlGnlIJnxd3uybFbUz
Bqr5z9KYR7hOUiNc8nwyDPIHtVuemq5FU9hxlTnF3DBLFXhWVMlSTTaJNUaJp2fSb0UFLkSzwkMx
SIrAVrUXetppFSg6L8Nw/q8d9gB+bYDUmmZOf/p8qiz2jskWp5HtMT3vMkF6jvndyMZwuJmR9yf5
U9cBf/GfEhKjltEGIG4RFXPPTwduR9IWGv7iuO6YsdE+jl8DlsQdQWbEcsy/L+1cs28BDIweoUYt
3oOM8J0wouFBMV12HZLXNRIAyhpLeRvtkCu8sj4exVx5Vy/F2zQoxLFUZGeHJkNQotNvWRXsIOQU
CG9Ucvj59wnOz5K4ltUou0/cltkt9YejSm7DRIgdVChYV7okwdPKiEgIZrzBUM7KMibhE46PaR4x
Vq2zWPHgPoEm2HOqxaZsbYB3/hn9GhVsTetyyeKt5t/fyPKhHomwSe9+Tt2GLKfwuoZXAfX/JXUf
B/zkCG8XB734wv667YBMSrhTO0+Y846xis8H0g7MU7oj+1Gne8Kd85hQ222ruNCtlvYZBLq7MhFY
hu65wziA+6n6M8RhmG0a2houlV/7MblCZXDr1dgYkGIPVcHIrFLmgTTxRaUR9vf7ni4HhWn4qjdF
uE5HaaQbM1jXMxlNOG8mr9SREBU5RRS+qM7lCIp6GmDzlq05KpNdSVUfM9O1wKHgeoLXzeSQLoyD
hzHJmI5uZpCHcQpVy0MVZ1wS/H/xe91Qd1s5OdTR68Pc6n9MTmQtm8xMUSbWtWX1oZCUIga4uyIN
sRX/f/e39UkYIBgCS11ah4P9N6JHFkOsRaAlCpFDOvcJHNzBgvY72v/eaBDHmyAH+NbYWrZCfQCf
hL89xMQV/D2J9hPf7YbX9S/1hwPV5rCzQ6ioPlRzCXz9w3vRs5xFwsfZmUoezwWsNOyRaFbYIAlW
Xr143Ng1rGuqCmWz/KQKgdW45tlrpx+RwQGn88slXXuFkLxD+NddEGN24pkZAHBQqzxZVUZurMKk
98qO82MvoKm18JocuvVW+7KFe5mASWd1NQeXBV/NJUNMUvKq1YbaIe3+ZQMzQl5Se3Vx9xKKfxMX
pddqeAkAcgK8HLDfsFmL2LTxpddSeewrJ3jLYYUDvwq+6EzpHuFanlA8UPbSXGF5a9KbEkfRelns
yE3MC13T220oGyFq1u3BYwEzKFlON/vHGaUSP+JBCDUpshasNlf1LMaFcdQOtQmHsccFFU8paM8H
PhKbnH1b6q9zXKkZJuK3eOuD/VfcVgEgXSmPrZ5zQUAeclQdWwm20hFiTBRS+YdDVn7Z51P9BaKj
QZfgyBbf/hQ0JptQwRQt4SBfc8GcIMXgcvgAHFaxgQZb8lO4lCqAG9omvCML+0RazcyoB/7Q4xHl
f3IRH5q0vloUrh7OHXQk64LgPSwo6JdEUt+26id0FDiaWRLiDYyEDbrKBLBdWudDVGo+t9ByBT3p
1OWxy4BhLQQAuXMJRVVlEeuu1EY+/3RSGSAwlAh7nUOeubQh8oIJcXpjBZFT7eaYJ4/xsS0yKt43
jmyEzfElsXgcOzXBa+DWAgTF2u2bXX6LHRp09owtBHmz/i43UiNnpCjU+uIXlgqF9yHe/HNwKvIa
2LB4z6EoIPA5oSfkuDZEDwYsXQlPhHCLieSONAnMkQwvUZW4JKAC8l6S645ry7MeBghK7W4AMNSv
fT+Izp2FJ85GS/kwTmxJvnHM9pI4c4b1jIBNDkvaoHXcAUh8g8/cdJwVzTr7OGz4FC9oP+y/WsCz
t4Hz4q1p8CK+/VejTnRSTYaLG21Y7A5Vr6+ic4EA9Ntp+rAh/nre7X61yH1jrm9ccVwj7K0+Cw+r
7c+IG1WVdh7T6F13Ofs4whJXZpYMydguesi6RMF644RsyM+vUOs2QBHDBwa1IeDrE3ze0R1cR4Zb
kQHLKheB6922VmkhIW1HgS5qnVzqUWpp3OUbvVLwlGQXhg5F6h0ahKVK5In7/Z1xaO+/59Xw524e
SR8vJtiGMGL5jtRP72nunx7CMKMBl1MbJZQ+CFzf1SSOv/yxRSCbwtxZhGmI06vJlqfa26we+nvt
pgqpT451ZIjimKX05rvszT1BC3C4H+tc3V5/xSRG6TGStoGiPtEX+LGwMlfExuj+krRWdvy0FUx+
mmJ0vRXsFzkOrBZFilsAgwLmv6kZJhaEfH8Z9Ei4KUwxHNmUvCYYrdvZUK5YQO7UDkamWOSpicXO
bKrnd2wWABqGqK0blnTO1ES3dbuTiDoBeEprlud6UtA4slcMN7lTZukfcz0fkCFdpA7hCjt41EmU
cim2XWHRGbtbdZI6UH6+CrGdubZEqOQ/m2Fr1lHFpDghOIbhCvsg6CdM50w6VCk1NsW9BGpLndfo
ihLi6B29UshjRjL3b0rfZZ1AI9o4MYS7/UvWQXNTuG1tT07b1skzjHA74LNJO5Y8bWtxfYcJKbVz
Wnm/vzbI8QQ/bDnXC2oMAU7it6Xu/t3fYLguPD3Cnw9lV0g2yf81L+FWqn7DNwkSh9jx3nA82WpA
I2iUrx55Nxl12Gwe24O6suupFobKqUe4c3pLV6N8RtIiwl4+vauOIs/s7AaOt8TLyJ/ZJ5nTh7tN
pTqaijG0GPSaiFlEIsagljzfpxqxmGba3jypu50NU5+lwTbh3LSmuB+pHjqBe0/IqObwAbVIfwAv
HTLjIf2ds2zKxj0a8C4u7biZa+hp4tnA/RklEPC+sm894hoSAvizL3z8jvwkdzWqOe5+uONAK3c6
LfaMMhXIgjCXvjssxV5NXmmWcdWftEDDZAyj2votNGqsdlLHHq65/Xv7WvwjDq5PYE6inhF1vFFA
NMh+eFhSwerjsMsn4mO4RmpCKK6A6HtlT91/HCqwHZs3j8uQj3SRgs3fV5Yr8L+fV0HQJ5Q1tNR1
jtA/BnsqQK1xB4lBWJP73Wc8FouUMC7fwVBUAvxGbk5DGmnlcG5UmvFYDai+kabU6RCD5Q5lFVgh
YtWBdMpkFzdO419jx2Y8/qcD37r+mRs8VVoCe/FceKpr10iIJK+BB9uF0B6GI9n3Kn//e/ZPbAZ2
gLhobxAAUqoC62HYm1guX+ma45W68DuuczYUMvvjYM/DeA2GHdBZxPLZ4lrAPwf1hLNv0UEmKQH6
tA/kVwQDWOdJlfAV+AQBaWFQpEI/FeA+VwQCDQjFgGP8S5jkAPyP+6PMnwpC/9YRahs6rEMt8y0I
4umqeGvxEXmNVjy8sIHHEOhLOJ2fUBXxhm5uLPQqs+dlBbjBOqDAniSqbBdXTajhy49ccD5bPVG8
T8m63RVp8ZnpyuiRdYXDmpU5GVCH6ctgTnIvzpLMuTfY31QxmDzOvwmG3nEmkWB25UOEY6lLV42S
hK7nqHxdlaql/jRyclGzBRIS8iphQIPqpNh3pWHwmn1viSdHi3KZLKG0QkptshLWsmH7dnuVt0yO
fzx1QhCrCKAzjN5/0fQYD/YXGoWcSzaJyTXtVf+NmzsR0QiEf0dd99YVk7G/u0mNZJbzn1HrHWvl
2RF/48FCcNj8nqXkpYAS0Po9FgQS1EkK9G3N42+kXJZRM5S4njkA610u/IJ+jPYtwvaHiGXbuB+4
pc2hypGc0SxUsIIQlzLUywFNx1GUblB1M4Chg1cle8wB2w4E1ksqJ4fgDJ/YGq/79cH20djNRl3W
5xpcruar3NH0pjL9rJhIClh28eSK5cF4fXq0sCzcbOIS5JzRJsUSZ/Nlps7jcaDNNEh8Tr23+iMM
Ig6iEaEnJpx+4UvkB30EK0lLdy5j8T5j9q1X8aUNGlC0GC26q5sf5Ta8+ImkooII/tNQ5a4GJjRb
O083PxmQaH86Kr2e1pDbPMfmyAKHl2XsQ2839JFakyK/cXb9JNcyqqXnAjKUTCYZZaW1sNTbVG0T
eY/6rVjsCQwb0qHK/6xcwiZLTg1O7R4A050yAlXmSonjo5FEcOz8iXjHv2v6WQJ6Yok1LF+zcd2M
eYSFJp+VsM2fncqyKsgc+vZ4agQiIFkytnjHn1g0IojYxfMnFE3nJ42ybw09qVqf5Sx9pzFl4rsL
peCtdcdJa9UZ/NCnS+42BdOOAv3uZnlyjT5Ss50hcHmOBf7SjqtAdJt/iEdqZ/vImtqnNYCfL1ej
PLseJNlOLTXie2OhfAeyc8AvyJFESn15A+ScH4z0wjy/qtPTq0LiIcCnO+M93JzXlbYIm2RC1Fea
ypRLt80eiajbRMdhP7WCkoET9XT/w1kbIIyPjHO3PkIFGW3TK2rr7UgDNDiA236tK0BGoBtBq0Qr
TO0Z9fSkTpLXYoEEfxLUmnm5Mxwj+b8JLjxsmObskhBiJCGnZ512AjotL+dz8I7g2X9MAbwG29Cl
wqWyKC/Ourgcv9J8FXJPpi28y76d2kU7P4U6PzyuHggEv2Xn0C2EVRqPKngVZVMvgUbe/1N3x390
m+fDrCep//Gi2ChqLYyKG56sZ5a+Hls1v0LuukecoHPVB8V6q5Kasl+5pjMBavQlAy0LKayzD8FR
XoL6KNHR+1/+WRL8vdmKoLR2L9FRgt3AS+566/yRt0eip3Gat5XTuQGn8qsXEh0CBSrQeEaJ2LCN
IrOwUImc+4oGs6qOMRCAIfhZvv0R3xMkuVMwLH7HH0UUIqABnMbHlrzuSYr4u8pDN9KGSA5OJwkT
g6ga+WPYKQPuppfqeMg0MMAzj5mZZQn2HIPvIZtLHnNoALoZJlRw9lq6pF+buQk7SxQaXdrS4Eil
xS/PuktgaixAo+O05GCr8DF+qxXi0k0D3TOe9pGSgravyrH9ygIjU7zKM787cQGbdFLeri7/eVbq
WTPQK7hs/Jo1MGSUi47Szqq04184Dfn3DfF83xN+ZKz3FbZCEAmT31lqFRQaUalgO9ksJzdo6NDZ
gx5lLVzoDNBMg0CAN2fa9CD4iMpZ0+lD4A6fpU4H5Ee3yMf/2wJFsmNd5x8GwFiXDp/1tB7ge+NS
fOeDb25aKfQ8C3CHCm62uLYkfYhCOjqoxCfegPxI0d7tqz35Zn5yLOK5d3LRP7WydqHcH76Quk70
W/2naSSK7cExZx+InlsBqXL7Lt9XbjAby4JQyrbs4eCIZ6EtgbkjnOiVVl56FLSGwWkJlXix+c96
tbqnxl3XQjJ0oz8fTP7ZpLAtny/uLJJmA4nIDjUdMQKGAXp2/eG1OetmbN3B64O4uGcv/rFAJMuk
K38CQYUsaMAankmjmFUTOZ5i6WrOLSyhzi1vdYvFG/pZBmhoge4aHsUCZqBkJngIKPkfS9qTF3VG
rcW+ZSAWbhIFAieDWrbGTzQ/R3wPYDH1pGkCg6CZR5Qga3Wde7yBWQhsLotiuTm0fbeQWpbe1Pqw
yIfUX92wRhGzSXxYWOFGNQJBoR99DQwO/JgAODb9LGHr6oruhwIGGleiBD0/mGUX5y6NqIcLB+q+
HipCQYTdgR4XA1DVdBqJjCuuR3Al1a9vkZFDv03NG36FsNpjDZYou8PcE7z7+lfexC03F9hTIYeE
ylAaaYwbbAIQamEKX2+SpSPcmHTj1s40073KSKbddljKGKdTpO2oeXbYpoOPU9MTZ9XjgPzrrI06
CEdBU1zf8XeLnQHzTiCcvGvtLE4FpnREdM/UMLScoxzEZf3AAPQWaHWTTp9cxBjnX3e5FFLvmB6N
mAiIPxx9lk5oCK056PAXswXW6sei0gyTsT43NQ/Oi9vioU3PrRCclaC2+OS8iJVs4cUKyXEu/uIJ
gqHiFIeVBX87R7WK2riDhCgbttnzQl7zQzkuboMrcutFD0twB2TR7aB/5d/vsBQ5SwqefV3QmWsk
eJQv6Kmgariei+z5JXhYgTDRWynuwmBbcjDWZ8EG/neOIvZRLdorK/gNZOYcLGgUugKF+55Uks2f
DK1Qgp8/tdgSu9aFhANW7MM/ye9uwu/oqN+DjXWqQ2BKINawac7maIwb/IlR6ccc3CNx7ltFD2Eu
lN15vyjD1y7bhCmNvEpt9eue5NU09phCLKwGgNYG86NHX66ACzs7qMtlKWafvVnv3LYSdnDLPpfb
j8KbdVgmQz0HNbZ2DBIyFbW4ULPE5l4yofxUGTnvZvMu/cFc7/NLnJwm+Zkv3Armq2KblX8qtvw+
9Oi2PY1bfd5xHpm65goEiOTuqgiIRYTKt/fo+nCshOwUT77V3pgXWB4LtReq1THyErQACqIyN0IS
HMFi7UK0cmNkcWLrzFM+Gbo45CwzuhOWi2AukIRUUJ24LJelOjfpee7pa//zPUggCEHajCIQN0pJ
VMmdD7gexSloe0ZnRmQxdXv3GOuiTmBTS+vy64/UarfKWKbn2dhm68aCUUW6SDjcCIInundbneGR
tqKo4s+EtJ7NPtHHXfUZonBFDfwf/zV25k4BwxX3pvJJYbzo+JUAYNteKuNH8sOyE6Vx7XjlT1fz
7ePOxdSYuqXSfTD2637rv/hqh+fTI5/cBuz+/Iu1qLRjDxNzBlOJs/dEeTyHdl+GoSzD+ExifGy5
YhrPO5jIvgGkSc6Ov3ec4cU4WIZIIGnLDJbT+ocxbtDHIwYBmav6M0ltdsQyxSX+5VtG75zRPIUe
hDZFfDORflucrkwx973dXMvPKVYEDQHsImcCzWTnnb8MwN6jTWgMN/jA6ENjQ9bedNfqYFJtoXcu
TNCycEaiLoVFc9bZa8MYFSzVvl3d/wIySnLbecYh99ad44w5j1gA///h20fls3MY0ckZ1trObdOC
2SUeBTmTzo0FlRiIIAfew2XKk1GJNhBeQL3YxK91+rdfv74jxFNv/LAr/3kFzXfgcQMNiRB+qm3W
Dj5nikKHxA7StrG/SfemZZOCmMQOUVThtGWTa9HiUbkX4sigAbRjWszKYGfGJ2EwaA4VlCLj2hDP
8xAJR0QFdDf10YOyzSV2c6hs1OVSkTnw4z9BTsoh2NWEU9Bv4AcnNiQMPFGNv9ChwZRFZrRzZUwM
078crMuaQpzcnlAJgxRgUXm70sQhbeO+D3BzXBOVZAl3mrXQUVLmTqG1eozNexYG6mlglGeGKoNq
Nvlneg5Fg2L3NXoLxtEQOkg64Zr3AIw9r4Am9x5w/2TbGDad8Y5Mx+iLzazjqL5LxwWZm6lX69G9
4+NxiDYEob8ugmduzPikmUknZUTPwZDxQ2XgNd95TSf0kXR7yAqNUwz7TaJWtyQ+IAAJlPIL/xyH
Bi8w5Om90Fa34kPHKpZv7PxLvOPSBRGGjdkbKLJqxT+Q95w8CoSd3OCiLCb/emp8E7Z+XPSkI48n
FkL1sBS83eRniWgouL5YC9lTXQFlBcLCjBF2+W1kFHNceGBFhkUrh2PzpXGSNfJs23QKipct4RGQ
5la4VE7eztA3ubmfIXpmB78d+5FX1GhkFBhKOVvGYAK5P7cqKP5MdlJlrSMUv1BPV/wzE2WdoKym
HJxb5Ok4VphGve2rDsMevtkldzzcp4Z1E5iSttWRTTcASjdwut1Ev7lE7MbyizhXvRrq3kk4VEOL
YKIHNOLB0l51mQLHa98wto7z9M2AdhkcW2h6fNToma3d+katmgDZ+ryJd1ZIIZw6N4LQNxbZy0jW
xQP/K3al0NPPEnCOL/dxucb16sWOQA/tGo3xdKL7yRj4teew3ks/u4O28rMaJSzhHmQnkfuBvOuS
f55OxIJWgCmtWU++3mkEKvdNMPVHSXKRUq67BvxzSGga0HkGvo2wU4G2efoHwCmQHDm7odNdoARC
2BnZHNYwogIf6zV6W3yl0RpQYAScaWPut+Tq2wG01WoEXEhTX/SzhcExugTEtk7sBPXv36MdvSSg
rBwIy+adO16bEsCCoc2TwXEorscXHDALqnbtRPHf6UozGXxwod1IoqtJafHs2C10pJSqwzcrGPVa
atBVblBEllLZ8qaQ5FPaQX7QNzJ4UjneFybDyBTnoeuG9VCmWB3yJ7r69KvsdxFvt03UVV9zr1Tx
gaI48QK1sFLChErGFykvk6u+yoYE8tEFlKQ+C4bXNIZ5ryb4LLaxoEmQyFAdondyT0mkK/zTba+X
GV3mATYldYZG+IqiUmbFQXvHQVXnn+70QmfaZMo4TbsCxKahHyR0/6Zr7j15w8/mfJbAGIm9+zuv
sPGlPoR42uKLT4MqX8DiyZpYhDLIsyKiBUcvOzUxRGWIw7PPPtbP57KaN31/TfmXsNq2bidjR1m1
k5cF8nK8XEj19NKZJ8df0XYUBRaPPmIqd9zLJ1Y0DjrgOeTPcfDlUwwZbn2krDW+Z5THtyrC4V0z
Kc8FuAyhsoJ1LENaiKjI6P21zbmzcvBqvGOAprkByjZTZnCMf1gws3kLN4EUraEpJC8cDfyAbWgt
5lT7WU9MBoqqqMmx1d2SPzOd8eXtZVPmTRh4tK+IXX9xrVDnMKXAVPQeyYopXK5BvKZW3j28pheh
4FoNgOi4j7iW0LkJYi1TZglSrwJI6s5sgvW0hJjLBhviZnIXQrwwfcyCmzWLm6vYH1X3IGyKD32m
yxFz6ue91Odkk/QISaoROYJv719PsHgNTX/xGORK/BLizMhtDJn/6nDuG2zgrlkTkq0SaaFiRXC2
8+CrSsnCAIVC+gUazX4MuIn0fIxrsO0PynIa+xWmi4px4yEpASLDL+/sGuMDsDiemoW1YfD9aMa6
6uzFGe/9Kz4daImqRdbf8wXs821XdEP6hx+eI67RMMHQZQBVzrrfXttiLmxmgxyEsnousIQ+lp7K
/FXfoGLXOEH3h+h7eS8TzLE9YdbaXSBXPoBAEk07NSss/dBlhmK/zqrPQCT1+37QsGpsfWcanD31
FASnhUQC0Rp4Ah0ml8ceeO0mzBCZB8fse+rF1MXkKQmiMqcdC6sIVUh0W9SE9vzn57PRGCy5BE/u
lYXjtqxeqBm5/RYFJEFBNMnlJ3rIpT1tkYAziDAkFcquw6+9qSNcIG9/CrYD3CfE3kqrzNCIJIlX
C10V2lpjydSH9D1Wh789gUNHCXl1JofqtxSOTkjcu+Qd5ChVT3NKU5a5nmHj7tpzO7C2WJANi7Qh
ueTfrV/NtusU5Uvd9FCxBT94H1A/uxiBer29HC/6akvy0rWeaenKRQtLuQ+tAAZWpGMsYaMedE6L
I4NexlFngCPDzbS5eEkYlRYS+lmfeZ3UO4JXoKfUnFiRIcI/ORVM7P3TfRo3elC3IQuiHgFSa/eD
Jj832zIG//10w7g5AL4wDafI0hxzeLwO0AmyzngdQ6N1YAfALCdAAWzEZlFqWYqgtN7RMp07CoYp
2YfF7Q1yHu6SWSUQMWxBcoCn3bngFbU88aHZbLJMmwgn7g26gUSTyahf2WstjPPr2RvXUd60vVXx
AYDjLzbdd9meIUak1StPgZd4yt3os+KQ2O2mvqZm+M4RZ2wDmlrPKZAXdC6B6znPmWQnOUBN6xc3
CQfsrfMYkOgWf33wGAJRw9sF29s7sWU7ksUc04h0IoZJp6vElqU4WeTcZRvJw1+csNVcLzNnXWLA
y7/l+ePdY05BhpWoNLmX/fZv07oKLvuokNCw66fKw1KNeBMbd9JaeXlxQMqMBmglDWYTIsA9Qlh9
v90DLYJJMfIPm+jrY72tk0ZkumSwebpc42xTfHJuBdzdnjf8qBWH8+c55V3Y6XT6DmCN/VKZ56dN
xprcXw9IRjTvHgTL9wWfDDPD8OUSn/SRQEk/MpMrMIfk55zFRu1AgOxv0y3CJ24EDPfkzWrv0b3+
hUUKfwOnVFCPWYDZ95pXiVcKmo10HEcr3jDvHZ5yjoxgWFr96bEfT9cDTE+lRMtOZ2Jlk9rq4F+3
ssra2rQeu7u8FyywXUnitsdCEnC0y1plG9OGFSv7qCDAlbIBxlufcVPXPZQvUQGsivSafe8semCS
XWP1NHc9tVJnwiyoqPDK4MVsp9K3Rf4tvs2noV3pzGUmOy1809JwIV7jJna1sP4Qec9Rjg4dWp5f
Uv5LXBjSFn5C07szfi9kjU3oSmziNcaSJ489J8V06IfXJhWueuugDWbomTQeP1aFhTr94mQVjWAg
AeWZTW00JlKoQ8TIAJG1oo+pX/pIIR8YdJ6pjDqV18N5qpX2XY925YYSJgsHtKYYO78BScAwqnON
9hotkfx7w/rUos5RiNAxQ2RTg3H404juSn+oLuP0Okpr/jdRyEGEyXZ2Z6/xmp1cQPm28P4fXvyn
4SHV7zOg+t7G9NSSVbWRbU5jRq4pEbZy+2xxRaQvNezmbHpHzNdFBg69RS3INIyde3Jb5FKmTfD5
0PgIlITAp4WVIeBO03QH9/YqlM2XVck3BT+CWIJ9W/9mjKjEOIkToUFjQDYMnC58dGVx1/tPDuwE
Z4XEV/sUaDC4TmUuWBZJNXag4DR1j01FmsoprHD8wxpXGEFcZIrprD8CH2NebIxVmsFoC3lOz2Cm
+8TYnaQaWKh5OSbcbTd8VxNVG1Y4fGTZ8U381/3aNnsCPIoYTfqINznKBveeri1zcif2GxFJWmIk
ZDGG4bLmhHm2Yo2+FWYYhQ0cldJw/day/ktwgWqH4Q4FkmpTmbbpOhQYd4nZkPLIUCExpzpa6OTm
UXvU9onp9ZjO4MzEVJMLXLxDfBTUsMS2Cd9ptZLsWtF90cvs27knDkw2DWjw5Bm2tbNXpKp7Y3fO
VgTk+oo0ygB/YmBri8KLH8SNPcr+5I3YwNzgyBlwhhTPPYvczjtWOUQ5Ob2niUERlmGeiKa7hfdq
rKUMluZt5D3dv9kaVzSEyTgrQ2gYAbCbsRU6brS9COc6Fe2xBOK4dHRvi6Su92Bp8hdftzvNbHGS
FjofqdhDhGU4UfZUjpPH2LAEiH5RaaP22k2eemUybNWlPTRAe9VEnzKWyLn7RUj94r6guBMLTwQb
vD6t5U9HVbS0iHeXDisU31pjrEdssKtkTsD4J4GaVSoQ6S8v1J49VpouVsRaF5OUZkzjli0XCRMH
jIyuFO0joX1pwOOLoEnzg5mb07kxPGCaSlbfw8oXwdou4Bg6YkptcjSnoFcIz4UKWyTEKI7Ki+ep
6wmOMBs5gT81CynvHWI8W0wzn9x68TrlktEMKPv2FHGu7PGFlvBDa83EHN1T+uNSxr5mx3PCxeS7
gl1uBbHIefqzETmesTbeoNduw3G+hA/s2BR687de63xw+t6qL9AWNGLWNktozGhhU8D8X2KtndRX
/3HJA+X24nVPqs5ZwRoOm8LZUBNg5D+tnwRxqsj28hppNgZUeEOUzXVkHPk6Lw+3oKk0EloiU8a6
bqwBVT2VNxMqqy/yKoFgt0n3tLqbvzFCiPh2HyoRIMHmyKv9UYE6XmevdYbk6KuZ1ILe9zxwLdlx
zER/Cey4CU6kX1jvWFFPEJBrdr38+IaUhXKjCFpnSMtoN91n+fy3CMN9FF8bel1jBipEcQEeRebV
5wWxMgR/0QSmEmgkfBfOPRW8oYwI7t+vqPuYHcGq0QPSGwFIa8xyxKUvAfMQT57B6S8Fo5Zs+sz7
VNnx7BYiwGUcNdik3QU8JgxR1/s2v9ul+ZjyvR9hU6tmo2VJwYxbSZRGoQUorgPCMmPZlXdLZ0Vl
KnmSVwrs7C293Qd18t+MRXSSzmVzPqaHZtFrhXMiTCHYLkZ5RI0JQ6f4j2nrF2yyGqLkslgeTPgi
wLXof612MeqUHDYuHPJA3Iw+88vKOhTg6Zh3T8HM/hdnHtlPYr5RvHAGqXeVXXp8vTb4e8a6Xt2O
jW1q0HqCv69eaOQfzdMU9AJeK+8zDVmJ45SRsQwUc2N/r8kVplOmOYGiD8gS4b1QhJ9QbcqnYrxo
hP01PPTc0EgbKUtjfbdwEtfpk3Y9Ok+5eacFCfYajXgwJ7oOLmAR5o5Sn9lbn3ciDOwnKzD3o8+c
EjufyaPk5rBu7rs+sS/LJixK7YpfLEcA8hsOGCi7mJtoSZ71b0sLu1fjQqzAUT43fJDNUGDR2/H8
WubE5hvJqFmSeMEWMqaRnXKOoCvgCQ2V2vturyja9Invbs9U5eLSsr/daI+mf+rFHcPu6GxoZQI7
5sEXo/aT6fQB28Ith3M3+cG38XgpDdn6zG7aCsO9SECmHnBrj3N1+mn90N+c0FuQpcqf0PD6TIFZ
DeH6NLG72Eq3AWNbb+ip/gqk1F/aV4EX19eiyp3OXNoB7HEBRQZDx4D9Bq3ksX3oyhxRcUEP/hDZ
A6EWmq0LEiRjzXqjWL81u2iqiT+9XCT5h81dHaDQrWbA7KecoEiTRSL7xMJyi2PZt03VNtqrF9E+
/8QEDfwRSSIIAyKbcgwDsIGhopT/ZnGwZtSE6jpQnwHUmpaJ8IKt8C4pD27RqYRN3nHMUPp+5iA7
kPJ0cyAXpDTCNUGGxJyrwEcFK0dP6a1IM4yi28hmuuzFAxmqfhnYGBXevySw7aHunEm1epq418AA
CYhRkvPdfLc3VPbyQxOIqv2XHr/dZyvA8BQgLmE+pkQFUXMd4Tgv50x89nlxgTzAj0HErkzA467L
M3+sBpHtJcLl0/7CL7L3tq5EOi66qJWZ7BTYxMhV3lgJ7a3y5uSJa7LzkNlXO2Ytu1x3NM2msvQO
cH66/b9bl/iVtj6Rsh/byYWxHjhLa3ifUI8jgU3dTLujpW4FOKGbRbp2fbEMLk0SbYfbH+EnBkce
CZzOAfxvcGBvWjEnF/2yNHC2Rtv3BuCA7hZ6EVoBqK/hpDv2SjY+iGA3GDzlthackenFQD5cGyS/
WZUtp4l49Q3ith/UVTwfLCcLSoAhngijAvvsoYDVwsHfmbisnLctH7fGyf4JdmCmgp6YkDr0GzdO
8+GZb/3LSIK96y4KubVyHqx3JpoEraw51+QVRMJS4XM9IlGfvsr6BvmgELU3w95CtMoeO4GHTzbe
paDqXpWJoCnKbblv9ildiQRd/w77h8iUPfGBKNrQA9lyX9ND5VrVktNmEa00Dr5U/gNl52PI0SNA
C5FMNsnKSW91issaTr/luazuk8Wj1VTYYiwBYPOzoNnDo18MRChuN21ClbKCoLV87QlcK0Eag4M+
xFco0P8a1XlM9APuHxhqWkz/0bhenhOz6U5VcIP/h/vss5zRNuw521HNIoVYrViQB6C2y17AMvV1
hVV5XPPs4kom80C3f3SS1SNwEzJ3CrIzTe0Bs41YFd9tCegz2jrcHjfYfqBKybmj2k0mHE1463+w
ZmSAHMTnFUyZyKL2ANqHo+zhI2OrWwDpbs/TjfIEKAKq3KB6/D8cd93HMxbxHehfOH8KWD5Bw38Q
7c/U9lhBJfTqx8wV/wYk2JuXS/wbvqZPl3SVAEaEPEhRS/7tDfvOqwLEkYU+RBHJ9MKNLBnI2oTo
xmzAosaXTcILyVH+WupYkPpikjL5e7I0ivcDL4FN+Om3EEMfals99Cxl5we4hlO+2EuaOuv7/BhH
Vx6KrP9V0xOstCAqUepGw/FZIux1+SLgMO9voE3llNMmOVtssk03tKp+1qP0esUXAn6r1JQTbJMM
CtadGk67QMRRdgSDYFKRWAa5VWtP8GGgQiWEZbSE3cCrzFsVAnky/73Bpbc1h+jQwAvDtFtvVAO/
9TkSDHlgbxepwgzk913UXyOjqILDEEERLnefUignsWb96nqUZN3ysvzVy+JXygpWqxgKRcc2OH9C
tE7jy6aHsanv71g6xKtQ80PbPPK0dIqrIlWteqxUD81oK+CBbLa/whZYU65l3vAgzAYB8VHcpzqU
HGKUcfdrbCPfCDBClBTNaXEBWRbueqG29oje+KoQ9AvMvV7jfHDVShqtmdGCBoI977YwGC1xzwgK
sphQhKzdCmp7ZE81puYZMdphMKOk4JVJ9A+wDjdSZA59cfROXNm32ymiKPsNDCaoBlY4IHUawhNz
MNwOfRdVQXNLj+k10qfRm163icZ7x1ZqQlPmP/uOxOJwnZJrHka2B7QtO6BLBb/w2G1asrHkEdoa
diykOQjr7mes4QJUcD9pBOlT1LJ2LpszocIXPyL7i3hPBvgHWM5lzyr27eLUuY9XlkUw4/5F8cKo
YZHhCbT1gtGg1Cap1eYgDy00zJlDdtssoGRwgW/XKrGtsTHDQSCgsRt5EicMRGF42/oy8Z0n6azu
TrfEB6xP5mdCvRbZQcsrN1ZfiLSlI82qPPG43PDwmXRMRfF+n4/PY+7aIWDzJi7AlAeQ4cPHqHdQ
JMMptjck0m6j4cgLyqkQ/2hwfjusqmafU2xcBxU594QLtJvgSYZmbZgU+dsZn1pkNacl4rUgVEtG
oZ8PYUOMlNZCK8yoCrayArv2gF+KiwfvyrXfVhYlAg4tfQMJE3OdTn2niImswmrSL6+QvYmYj3oO
uSJ8Fz8U9tZa/R3wvhYMtNkFxHPrRpl9h5WJGqJeLFMCSfHRWc2De8nE4PYej0KuCcAmIOlMdesU
fUzqPPVzURG3peDE++GjLJetD2lA+9JSIrnF9GadETiaYDm5znSg9FR3NysqZPTfvRpBVJeX/BD7
SaoEYeVdFcgV4mj0yyu/GYefkM3+B01VbQSvKDpGmoEfAAvZghsQIN9G0w69bMDovmUcT0AquGxE
ow1oruhw4+aR94l2bAZpILIjyQUXJzSIycSRVN40qvYoL/YTG50ipWqJ619Rwl4Ne3A1/8khawaG
2ul8NCTNrggsX2uW3Yd3BqGpqRJrmq69juFO1vXsYNt5EN8fXmXwto7FJ/iZQm3gK0cy6f7NhmWV
1pSy2q+y/CbrQ6Y9Ic88juybiGY7RVCsQ+q/feIU7/1gCZze7BUIj7mgs6wFoWlQJlLbEAE2ggm5
W0q9ktxqUKL2o6oShtOHKWIeLV9I0CynFcp2YpgqFLEpmyI5Mz38BWj0jccI3e8iLsljVD1OKK6Y
A/N8aD4OD5H3n58GLNwy4ITGnAQYmKdLO5SDujea6f4YVu+5+V5kBpLNuCR1ouj10yqMP2nkfWH6
0Mqtj5jEe2DwXGsX7F1H3K7Y8sofZLs3ZxlJtLIw2+U2BHfAb8OMeBbE6j0FiAeHp3vn/12zgHjA
Cp7wT+nbtkg81gwxeWGsuC1L52wiyRgtuh4tksooSxUKoTDlPsqSny/JDC1+3AOFhB8gbPCNSUen
HBg+HxhYuDWsV44wiqGjEw4Y5jdB5/U+sSHfB+5Hh8umo/4QcsgztWT2OfDsMRdh53ZYhKW8rxGx
7bgxglPEhjvNRoCgaFyhpyHnyx7SqHka9U+LSJ9dPw28sJiBRziY93qBFnkfcL1AZHwbvMsjenq+
G/bKFY9AANM9JPzcJXMOt2CoVapJJheh4ATO2QPRrWeDtQXuu5AlgdLq9SQPxTLtVYlm1lg2jkbp
rlKGdY6MnZL+knqnPQpeY3jNjDxBq0xU5AZAOsXjZoM+aTjTxaAoYAQq92dgpeXGauQagpL2v9Oc
IRL4SbUvnAgOWqKsYmNGHhjGF+MI7pGpjFYUJ58Z2bGHbTRvLsrODfqtshw1SoLDp9Sui5TFec0S
ObcXCMGEZOaB2oM/VDyZbUyaWKoLgHmxkBGH86UtxsrNmFqOetCJgMyHDJZZ6fuiEu8Xm2G2mw4j
yKwK9WKObktxJM1kIUzdaUxRkDhea83NAh0y1HFoc4ug3L0M+JmXAn0kkVLxpyUd6mDyNHRRdCVl
Ym1NBms33Ld28MgIXPtmWXELy9IwqBh026VPqrvcjnHIFX0i9vDkZJjijCJZvR/trUh20dIVqSSH
alx+3k6lodl6hhaW02YvavS2gEqd8MgWvwrnoWF5+9xkPGTzBROWKO2AOKrddwtKDfciRFAOWd7O
Vk/rXnISyiYLRwPCJA48piMuYTt4jD14UX7szpn3v48PQ1zfK7uqJNT+6QSw0M5PWqGaH8pbQTb7
aZBTk2Ex0l1Uyl4b6Tjr0k1qFnMb2Q2yVMd6hPTdvO6QJW/K9eQq+jVkksTRWxRATO2BKSHtp27S
qbXZAwtd2hvh3o+PO9LTnODvqHnpRJbUmE5F1IV1ONc1ALa6jKbu8b8uZlhvO4/JoHswKd32wqJV
vdXKP/hV9u2ori8z1QA2OCOIdqJZ6z9OeBMTaqz74vTTYKcUlzTC/v7hilqwYU3BOb4Zp3eEGpWW
SCqE5QpbyCOve2JuUXIJQGLb7AYTNBVLzanMmPZb9kpOXRVUTyuU7qzMss0VqxmjD3GOI/wbgLUR
uiSzPQy7BElopGGBISczvHLXFJNIedr6Iw2jEKueiSnl5bS8V98h90BDj8hM9Ab1PLFHKzi9Vu9m
lLvqSl28jPiAiFeKxkFHfFjrBGlgf7at+Qi8N7bi8u0QbaD3ePfRkuQh8T9gKRYYNIy9vUJFyXn6
hWtuoEDTO83/wZQRUx8qViP0mcGSNasmNya6TG9LBaEmSEFYgFDG5JQYHsDwxt8Z+ybVCWHjbyKi
FDJErE7YQrlNp2SuznaeIxmWqDtlpsRdNtm7wC5jVhUZv2Z6vDjJb0no3vM4cNgOm0O+sGO9ie3K
APri7AgLtrkcXjgAyfcjki3vgTXJrpkMf4lgH+2Qx9tcdNl+U6svLJv7fdKEhhUENmZXg6W0gZfi
gAmSgDOdx2RBEZxtyi8juGH6hNFxZR2AyM9s4P90SiDRX9SC9pIwblq0VO1bvg+i1AlBjDQdKGoC
AX7qYwSj0N65/hnTJt8HCL1wkYL5L6hk6Aim9Sm8v4DThz6eRwLH1Ybfu9iEssKMPQMzUqckhYH1
39sJy6G+NJdgyvCk9FWKz5IZXwez23SF0nV2ZsfnYgcLak+8BZ0t5iW9+6nm56MPjycRfBCnp5m5
zlB62iOReZO46ueaL69HtIbiSFoOXfQ7z4RwmzqvBzIHTQ/P0QwyoY0DL+fpBVKiSl0i+u73z/xk
P92wmzj/FV0idugLijvq0+G2E4+wMtCEKyupVzenY0b/PI3euGzI9WlMZDcU0UFaKtkA0i4vWfZU
eWNyllMDS93xxRaM8oRto62IY0ZqKezmS0wMv5zGWye5FmbDLCg4RQ19VU+kaIvKRJx5eObXz1vD
bwUY3qgWh5Fi9hyi5J2gJ2VMzDbk+gCqevRPmmfrNcOMbKxn88x5J4AQL3g4QOodAFIpk6mvk3AM
quAsXAPeAztrct0Jctki7tFRhNm7yBui/LDj9W07ug+8/jGjQg/WGlNpTsWYl8MU5C8dhmvch+ZK
kBauJZt6T8pW/t+Zerm/YigvRVlh5EpS5gR7I87s2yLuLcsM8f4iHZIMz3mcsSWQmPw+pbn/sMh5
FFSRpzuR10vFyZL5tRMfgsZu+rpp5uTgP5/Fxf2dIpEFTzuDEDwcFoBXPQ+eC09BG7GqT/w+b0Wg
2bdCQxr8U4DC98clQmZkJOTRXMRBiu7Vv/TmaqPJ+L/tamSFbxfLX8QUpIwyK8Fi5rPPqXuuVNey
4QXUuMgC5mVPOSp704dRepLznzXRfzhTQETRbffmFg0GpTMdT4+/AWQzrpcEERFNoZe/FokNyeyI
M1y3OBA1KzIvnW4qZ80aTOIQl0ypDs98izcBQvK64FaNyhsNKY0QJ3DlzDXJ8ik3UO8EKR5sFCck
xZFqDXm86kkk/8gKPqmnVKbzceWsOm2MBIBWwEY7wEBq7iTtqgcvusT3Mi3HREYzOxCNfe1835eK
jXEUUEBIh7c43tOy3mCDNzylmlKxemk5+tFv7JS4sLgAQPfUisg4s7tBnau5Wqs6BdAD3Qs5suGD
YWY1yvmi5Kcb3fa8CkEbMVokKeFrTr6up0j73A01qzBQ77TB77wZ5xgklRFWHTTZAeaHyhwr5bUF
jy8lXbQVv7SJ7UFSm/RDFTxrS1ztK+jZHYqF9iq3udSgt+kjdaxYHdu8N9RLB+W8QGC5UB9qyGMG
t70echVD24DzH1UJJhhG4enjPNbNAxqGvRhQGtXjbl7ANWep5b5Ksi+AH3XdxiVKDyOsEPpDq/2L
JMCECVwJU18QWyi4wVZQct/V2S4hGFFQ3QIA78IxkAZ8sp8NRdt8TdnlsdzVFWwXUSBm+VT74bWb
CA1hqPxqnH4RgLfyL6VCvDM9jK3ZbIhkFUT++BABcjNCAYBVXMisepcMr/zx82I5rDiWLA5aGgNj
ORsBYAt2K1lEPeLnB3aovUugHYAEq+XdQPHtZ6eqg3HPUUdhAwvKKjREzvS+OeTR30RbIS5pmMWB
tMP80LIpickdUGO3frz9YO+eOxxQKFpdNUSTS0ENsAVPHR5JQOZLsELnmjsiAXH3MPhUzteXmwl1
laCUt+e+RTFDVCoOoj6QwlfxRQJL1Uj2EKWDGxvYBqvbJafXPceX+FsFlydMfnhuqocs0Nn1gzbp
Hq7xMb3POk3Lb6PRw+T+xdOxqOP2yO6aONrxPLsIXK7Zdin37mLa+nLG+9gdA/ufxL4JCMU+nta/
IgckyRx7tjwTByt0IQM2ylT2m665KdM2+/lkAvaWV7dYSaLUGUeo2rC4RChGyX7HzTeAcM5M8fAt
8HLoxO0V/UP38UpJaUJlRglkNf78Uq0jT2urW4e8gJ7gH0NBuQ4IiWk6HST3TWg8BRdPiL3uQVyC
pUMzSZK44Xy59BqZ0kjpuE887JbOke/s7PcbgC18qrF2ra6AGkDqyX6R7m17mBJjFrSMXf0kLxY+
bsfUPMxiQR5FQ+Yr/7Fxs+80rQg3luKEDZ27qKqL6H2gyGtWplap0O2oCKipo9LK9A7/TRf0pdYe
YmjzhKZ4nw/Yr7U27fM42nNuux+IdsTt+ZZfTRO49HdQX4Ct3juhBPcUxSqK6rJuFHTh49ysIKh1
tCLpIFQHP4VsBZJDknvvxa/Km3rDqtzcv4Gz6PccPuLHaGgkl69lIt/wu0uvmZUE49Sg5D8uGhZn
9Fi0JTckLH5rqSqzGeDFwj0WjUdt1qD82RLZe7cEH5ZIc1tIVxs4yjrTOCd0xgn51huyG8iTkX/3
JPv3hMKzmKOx4BREMgwPHh4eP2nhaBqS/LNfzrf9/xE+B6FIaBnEWc1qvdIzQDKUiyf+TG4biwoa
qv8NvqH841wpbMkS9sPes0WfPLuFCttBqQPlDYAgLcQxr9NEZHFpHY8Y25/YeAe9gBoFKfXQaQoz
/LlDAdMt/jTk1m1EtV2x80Tj1m0ZGZE09E92tu9qB4hOFuwC6r7bQTT6Wi/mh17hAPx/tUPzszuW
EBHhoNI0ydWfFzdN2rX8waBCQ4nz+cGGZcFM55lGVXOV4pxLOwGuZindiy/wvoYZBcl8vAUMXDlF
QYNCIGegzXuigh29SNBLRZcf7k2UBWexH+XMwWRiGMw6trYTKgYcZIfbUwLH65gD3tatXFyuuQ+X
W0HHGhyIo4aqx36A+phe0owGFXWuBwnQpCelnej0kWNYIF3xPrr7FEb0NH/0PhvKjDCjwcBJtnOw
5H2LD6B9+HnuR9OAuRXinL/fZ+FEsmHb9BYPTUPXN/UP7WMVYQ/upbIVPwQrFefSNGSOkp5ew949
S8RgrFGaarSSEF8llmV4uFMPDs05yv8GijmTQWwX/WSuKrC6QTdGm5LNtSQEbUib68eZv1ORp+cm
uhN/3ks3OnOzRnGAA3+tO+oL8AcFq9WHtSWfvh4B/en1qbFCVpiLtRtDM5i4Cn4o+VS5stpe0GSj
V6oZltVezJSKIXJXskwxkuBEwnWCYNLpjxUI9p0EyQRgW1hDO6E2jtlKUib1pwrikkEY+AlLFd/P
WZcxxDCSfqpThtt3UXuJtErtL9btw9Nx+Ek+VojXLx5tEZvZGlbUBt1miEYl7KQ0j0x515zjlgcg
63ZYsNFBK9MFo14podEfaUu9S7izyVEEm8iTCeIyozb4YEsYlnZVoQXLIN7KGoRMRKHEjhX+vx3y
X5GtlpxvxxrgliwKwHgI7JJzxUgtkioTfOpTt4xNXBok6wHp/RThtwoayAL44PLL9822hX8sI//C
+Zbx/7F9ybjCUDNAaM3WBPnJSjj0zD6/Ij3dzO1F6woPhP/7ifcnPf0Mz3uRXXJvqbuD+iJzCeAF
3A8HRcGQiso56nkoqIQ9ChmuzbSy+VTQLL1Y6EI8bG4lb0iL6lxxvkecHrsm88KfpkvLu+PiVw0T
dZ8a9CVUausSzNjYRRa+RRFUME6c2YcK9O45yxLLLdFHC4AzJu16gmZ19bd7BKWfT4epMryDWUBd
T/KBvt20Dyg6d8hku0jdcpvJqpU9aVVXJpkOhcWhxSGUBKNn/LCuBkje6myxN+MATtt1l4WMghjb
FQWgie1QziAS79jurCIbruMOudK3OPeoccMWhgBi3y2yqztEqIDCb4SC1VDnFg22I7AhgSVQIqfk
Zn/+ucBSMJnG8aS0K0Poxtq5xrFPeTaQYbA05Ja7lk1C0VoIburZoVAZzvKOan84+TLSt52EsqpU
tTb9xJe5Vnwplamj6UfO+YwfMSTgGdsVrWCum6ZtR6XgmVyogp/NuMqfbW/c9CThwete6wTy9ydp
fLQSsfdvs9Wvzb8YQ//wJelogH65l1T0vegMNR+H4KIfnRwOtKZItGxTiuomIlVN74dvKcVFHAsj
WA2bopTs4CkgQuo6+PjSnoMwsvG0NmZI5YjpcfJD5lYsOaFfO/gQfyoejZ+0kxp+fZAEviUL4EFm
XMz8Ywo2d6n6s1Qm3PATvYHtq/7hAYFnm5A790SUbmIb0ErYvFjl/UHBCBnIgh/xkzLC59mqWqGp
17Cnj3tljhTDm34pKlU0PxETEzPRFbPLQJZUf1gtQ4EYON8X3aowbZT7hTno9GRHUWz/0crPdqr8
eNWHJ/jhC7shqP2iQPFMQ4AJ7a+Fx2g07lrd8PSaYU9Rt6lwgDqu3uoZuwCyy6UfB6yrbQ4Df05U
rYFRbw8RoY173bbMqqlgAnV3VY017MExLHYY5Z7MsCNjoyzghCp50qUmqyzZE4MBGPJk2CfkqIlg
FwmzUa993Wqx+KP2Open6c8hW7ZB2ZXOAoRvi0+zk5TNqYfdw28OCjAUgR8Dvk53XbRSnQC8ZSKl
P8Sfy3jGG4jyJCwHN0cHiLp7GXqait0/0qAQcNICzdkCWW4ozvA9QHv1JO07/aqKG+xvA6JTTzL6
SLKKZmcZWkZMxynB+hjcN7aU0EQYrDWFYWVnVn24npUr/aEOGtqBVZc/lDsHzEBD7+xEOGeuVD3+
7CxGYQao2qcBMEwRTZFqovI7UyvZLgpasR8m8T7ECA2KA/7WaBq/oibAbZCxC9U9GPrPo4qIHk2F
bbmSkPnfNIwc6s5CEfpYgDF7ZhydT0Eq/pw+uAmC6vSIZVrRCiCieolY/5lYt6H7PjfgvWUz15HN
/R4okKOuSFPX2FjiJBRrLpO/l5Yrj15dL4/cEkRoKYg6niMQ/l7Ld1qDAyUF7EZt2UVuZeMW3NE1
jYrO9Fm/2p/qv6seUCbI+MzMYZFD2uoeMZLCaFr47V41+ux7kV3rhK1EtgXNo2iXzBfxvaadZjut
KMLQrIabLozK+oFzF0/NijihWiz7Xs1At/8qbPMsjJNoRJyL5D87AFo5BMLe0x8okWGAYAyFqHeZ
f/+4qhy4eFsHJLwHUvMG/1jgBl3ecKfeeYQI/X1LRIgsa1bMP2hPniscoBcn1bdi0IorJsa0PtaV
Za58PKFc7fXMpd1bTn12aMoWMqGtpkz1Z4e0g7t0gF9RuJKb0dBeIHDGDv/HIEUOQFJLA+SpLZ0P
7vhvx4wqjQTsewyXxciEDUkIVExxk2ZuTciKmAHSqqALCYmF+mioARq+Fc3x8k+0SllfNZA8msNk
W+AcpV6gzRLaBh9caj0RhmzX2BbY0Eypp65M/QEFYKakIna0VN8f20lAEtjLNB3jADUFBIdhxKSz
MAe8olxIRfjsCtV8qAZGYWVIM60oCuNQhekCQ/H+9BDFxTi+eJ4poQpwSx5CXOi7mEAPjgW7H6cf
jfoLMdgEbzV6FeSlEW8aVoxqN2fGXMKkWFwsfDmqHb9Sf+MD5aQJ6/6Y2uYFA3+JiEThFH8+kP/2
0MZVwC9E1KHuhvr5CmxXRx/rzGyzjATutULykLU+y0RY+qY/NO4Fiw7sH0S8E2nlJr6LvdVBW73m
KaU9UoOLNPVNFWCcN4lYZL4u1o6MVlpwmyxgWvu+Qa52dUXZF9wxPe4/uJ/RaXAze3m1li3dydj7
x1owS7V1LVZrr1cXNtp7ki24L3cG6LTGW/PZAoWhlJUKAcBha0nt419u1KeMOef8Td84Gpsx5pOh
A13sGWjrqDe5+ZlYfRai7n3hsTk6YzqMCpYg2q5Yao2CrNzHrAK+wWGCbJW5N8Q9fi8RgVBSb0m/
bBEM9Yi41EZmS2yp9uBJXIutAZYLrSn2gS/EYbl/Pwgrt9rBuevZQvURqIqd3FlBHBaCPtZK4LK3
S+7HqiZ80JGXLcK2ssacvu0uQKxP2DdwWS73llKan2j2yYfJwgGctvu+H14Php6PIN+q3Yvy996w
JgY8OIYEgHWPMSqxTaB9JkxwmVPVb5YWCI/CqqOs7t1PMfoCMXd3FBaGVBAPcZP79o1cdv4TkuMq
ndaN8fCAejYiA7FfP4zsAr4p3J73L1Ekjuo+ja3b4AqWXTaNuh5BnZn95HfadcEPFuECYMgmvjiE
v0FcOIvzFdegvJCmXhDucYP0WlUM2gmD5Xg2kqvaGkJ7QwRJnZKL2PcvcsGLqMR9rIZaOj8GyfGQ
B5KgO3UrcJyd85BS2JQkuEMAvGfZPU9e32lM9AGopUTHza2Vxc/+ryuILxQUn61JYtYZTsnMresD
Vnlod3YqnbvV6cuFTJPQC2GaDVh4oX5mkM2eNIDYveTfT3uCvPSR+73dSHQZOgrRYBT15+bdS4rc
llfkAZyK38j5bm5DKEu6VhWbvJZV+zVJ4en/m4pqdwS2YX+aMOc4wOK7mkK+ZIYA32X6RrIlN5Nq
OhNyZ5q8vcxk3MvMBT/xSjwG+KrS7xtEqrAUQqgefAivJZ12EF+iwlvZClo4KNh2EpmYEVAnNhx6
oU1eEdqve0nvRYWC87dAMgFfwGcw+KjIUqM0AVaBk6aMyQC7deeuKk18dDap+iwRXMnYXFqfDi9e
P0nZ63dc0bXwpWZyJv8LlqGVdJ5NGZNi8D1qNvkd3gMSKhMJweGg+oTfzCNiAg/tYKIPaN1nyaKg
Atk+qGSos5XDnP2ON6zp0wNEA4SRN/soLATD+zz6ZGv9tfnETJFbjIOsjyQUs0JIt6aMmxopw1oh
DjHkSTGkG04ZOK0X7GxtrxRAAWt+L7EpRuXNsPlD+m2v+PYqzI2Iaf+7r9BMV5QjFWxc9uz1JBS7
+yjJY8dmwaUZwF/ppRoA1xj/+eaEKmq66BqjPloT6Ek63/pKLlhlmKMZnhCwJCJmBcs2cv3n4nRl
5mV7eKiRvNXDRtO7lPr7rlkbLKAX9Yc7zmd3FbuV+qbqXfjSJ//12yRiydaSQ1vJ+kzh39JbNM/s
6tYmrn64WKsriEyaBojuskKc7pYRbGwQShOfamHOeHejcMxf75qWG9edTME/Y816o+1cwmCrqo6e
bJuRfKBiadcT5nPNYxBtDR7z0Lj6oqxzed5beYlGzWpNvVbGr67KL0JD/yJOk+Kt+jw4AGeSncjj
Ho5eMJ9zyUeR5cRmaolXk1Z1yR/EVMLjECXMhYKx3t96y1vnw9o5mOKbSv/Z8wSoNyPZ6ug+QELl
FJ2XPL8naSCRCWrlctrYsCM2FzfyC5z2ajHF0ZZXZawmoK5wQdKrs1BE16xRifb+pFvpHzmHNJNW
t7+kuLFp6lFXqVF3zLCkeY1+wMipbCGSZTrIRnsq70olmqWfFKmIV3n7ktXpOJuJkG9K6/hn9X/B
VjJKaimwCT71o/2pgSQARysdwHHSPk4fA7wo9VgiiCqPH8a/hJcKosRsppk+89AZ6shcCe3gJpTK
aSb/ChqWScXbK7Fd7mtkwX6wwsUFL57cheqpBw/3PbExSu+ZhUvWFXy6Cy7vS1+oApYFoCZdH5zB
GCDxgbZg34H5pdQHO2Rm84JOrRU0MbFETFwXSBoxIaHqWhMWG2vf7G22W4IPW5QAUToXnuzUsMAO
YV4AAh+f8ZuOKD2EzPQaigALLhN3ru4JpRT+PHrPYfr09TmKVxtsy0v70QkoCCglLYhFJ5q7LuSy
JJ1QGK2pS/XwJ77m849ZtlikA3swXT7Qp3WOkTVGEVcWSXQmt76+kLx5ytXSd/tm+gDMiifJWJ4u
m1cb1RwyhNrAv7CZRvOKAFZgl3P0E5mSeunkdOxn0zPRr5Ytvp7+uIOSbX3jNEa71EnxqGDVWkiE
Kw/8+NFVDHXHw6Qq2Uw1ixIKulhM3LO8Tq+r9Bzpxnqz39PYkXWJpzQK4ClXt6+t9x8rezrmeBV0
HamxOnjzdepO9ZIpCf7YB+kR3q9MfNGtwXoq7LNFl0clzOghxo1qeoBqFsS/SAQUtaaSTOR51DP7
3q7bkw/2qUADauJKkUfcQFRCd9E52tVmgoC7c83zun6qcsK8K1M96DWSZE/1ijvjbP3VsqVEAkxR
HrWIHrLAJqOWf49RrTRzdoEGWqnZjIL6sP72G00iEDuLB/+Q9YSmHiehHDSWnmOb6z8KbHtojawL
3EsOaDi1GRfyEfj9U1YcO+z2k0JshGTVtrucVws9EcANgRL3W9Dus1NBkJi5KfMRt/EhQ1kzA1fa
hMrynh4jLLJBJV6n9Bvdrz4S5ixxLMXjhNAafZV1LUqPEsb3EaUriFgaWwt9E2X9dHT8jOpKo4p4
u+1DrYUxGJwKpOkh+2fRLEluwMBv5s1AZbAmpJyxcXcB0IQ7cFCRqSbW2cEs1th3MbqYxVw/9cZv
0iDCnmS4kHPLSWcR+lbAwa0oj8T4txgf9BT4dvIcGRgHRUOqTkIJK/ofeqJelrfLG1478wTP9/EG
S3nZMWfIyPPlKWfMBIQECs+6aDLVA6WFpEKvlWPk11hfnU/FWGJLsxsVZwjQxbMI2T4yY6mcFADM
FmPHnzv7XOtpyDOPWsntxxZfcFqFVuW0XolmYoQvUaGwRWGk+zyZJVgTi6jgZEvvnOSUnh0TLtwa
Fu9y/coDa00F86L+pYnD5igpgGuwHYwK2aq59hIZJYBPEH4QJvwEE+nXwjWRdKL9U/ZdTeJbz5Kz
RQhvqIbEqvdLUqEbxX+XVbm1TZ9awtBKKqvqmFMGAUftaZyvpSDvhDt3spuQsvTce3dhsI9Q51Ic
GMiiqKPQOVcL7rmIyE1bCPOHV5GN11uQGdh7g0cWVVaQqdkxghmiWrq7rHClCgEydDfZjLtct9l2
hOfHBGnggBv0BKtWkP/jTOc7c2jRGiKiAMxUdAmx9ltTQZfwKw6TlO62NfJsfVTuCmVLXzTuHRrD
qHLsEnZHkb6uncArVi4Wc+mIQN546xz1HzUxUoXT8dYp9jD/i6a/QIID9hxEl7IIWpFhnGSOmyo3
ZlHb/fEr2UKgt7+XHvp4lwtwAIn3uGhiiZhLqSBS8JgCcriXn7wLePx4H3ez08GayQdS4PgNoHXA
YK0AicNb+Zxb9a+hPeCW7Cqu9gjfdTLzNC2n+LYsefe+hftFX9dvcSmBVKJt4MXAK+TcJHsXC9JB
4KTiON90n7+wWqxGg7Zp9688xmfSBMUcbb9KW3WSad7uZdXqnJt3mlDeyxwrhcZbxmyKSp4KtGry
DjkqfDsJ9fCBpvNazK1NF7IDx5KefPz1sCCKtXqoj9P69uYYEJvIm8gNaBZFdcxGNnpbVHeSFZIP
3q/v47l5hWa4+yDgsI9uo2Y0M9yViyAWxX9N2sO2jFfxin/51Q/lQcFjxXQOHFztaE/uTglo6Qfp
cn9Vnib1NPhxg69d7HXzQds+H6sXM8h48RZbVatzvrgqfocMJzV9heZJYlZLzXztygn60do3Icbo
BBGkgDhY7qQNpEBdTUKNw3VckhNJKyn9hTswlvVAGURO83tXCnzIaAHk9Qeql+s/16TxWWhb8PSZ
AyGjFwV3dSOrS3yENuvbPOy5a1EaBJIbzvAL+zlH5es6TgMgEiJ4lNsHV7r6ICFby+Dt3wZj4oYO
cPz/91rfLBRjbOtwRfkqtKSAFNPziBtamyZMAPBcjzXjMjrHM0htV2ho2esFG8YR3T+ekQbBPcKt
NCMTbBbtsIWy/vp653+wjWCTyLZaM/Fk+PuygjjU+mP9Q9O4yi9Thblfl11btSqctUz/1Lg1HqjC
arPVDOyZgbFcGpRn7IIfTxqCefPK6atgIfPl1+yhGchRKzAuZa4lAvg9/re7jBAtN3A99jSX7vfz
O4NGO8TN08e01PrVvzCLzECYHNHtEZi0JUHDgq68yLzbHkN4hTH946/GnqmB5KdaFE3JzRY4DvB0
nWW14PcJpv+g4ezo51hZBZwyVRn3Gqw6MKU/l/9DvAumMuNDwzLRUZTzs/iMir9E3q153A/vFGEq
a7Zn5KdHD16ED5Fzpd4VSTar3q+9fz3JQ5O2gGpS2H9LGl9DP+1G4tvrCX1alZRz1Hw4CMuTH2Sp
0tCJ6HLdZMt381+KD7Qrrj7KiSrjSMUDnAr0A/iUcbo++I/JO2aBd2I2tlVA4U7b9yyQfkuDlTVC
gaeHUBIeFCSUbcusl3RUZkvkbcDDprKg0hdVz/nQQPbfbIFRuu4M0cSXwScaa8kHQrz+20Y+1KVG
Q9ezrOa095uNZ/bP7LM4Z0mkl1YL98vyKY51qfF3PjfsfTDHz3sW27C+3NruNLm6jknDm/UHpfEq
N2vLy7jQMWCwZ/TGs2JKZAyYy2koTOhanf+S9THgkMWdiF0MEy/RwbDEuJzwXXrFuwcMbxYgQjYV
hc2rCD6Uk/f2t5s8oaatpkROp0gUdW+OQuFdV2Zoxv+ArqKINRv3Y6ZS45Fen563kyULAxtTADRW
rvuY8LbYlr5IMd4RTZuu9ZsKDdux4GohwKfeqtE+6G0g8X1j6ptuCEnIeYUtBr4iZZGbYyi9WsRq
/Kp6HxorZeFjZtUbWQwdCVbEalqGriVq8p9hGyii7Fbw+ZboB3MC62/7+sN9KlyNB1PuSMoGHlPp
8mhOipQr3D9k1y3bXvmxAPugAKwKg/tEsLYbRxe1EwWuJZNtrQ0gfG40yoXuBl+bhTX8+jyQ1Lyx
rDN4UcaCJcoywJrPfsfoOnSA6cPbufTyUh6ZCQRb7h/0JO3xV8dkSQOmOTtEYvtPEVwyLNPBiypq
svJAX+OsV58h+kodI7P7sf4L1XyQrj1P8/Y4bHC9UciSHsDt8PnuSQEjHuk9+WCeSs81bD30y8DO
HtjVfuBvs132UXhO5Y4ijps6p14RfFy+rPlivFO6xWjsP02FShfkxtYbq+TisR0bDtzdwvJsu/ot
9ZpB12tQFZenJHOwYFOdJFZU8RKb4Q74lW4YlSK3YGFOuF/Xheu15MswXXm7IsIhWb3UdnLQu+0b
nju+Ji1b0YO5h8AcOv6Zgeheei0M1wCIfcLt5XKcV2xF7pW5Ajh4FblA4Ql8oueuiRAT+2Kfr0+r
mb4/W0498dVKSkrrTOR3F3pNxrdx7nsNMPjt8+qLayGBiaH1h64v+gvPZR6I2a0QlKSD7B1tFxxb
gagJVborH8GP5fJ9EViCOJXg+cRA5TrVL17CQr7iXDyP6O10HL8K9GTeTXwZwtEmKFxSd4Na77vs
H0HzDcPSd9hDy9R2p3hWsimTnWIT424Q5XUdyvxA82QDAj8I0vIeAIZq+p8n/fA/QdjxyQiu5xAr
m5h9mGHWAaOx0MbVQ32otxjpUf22oXlIDsAPd1x3B316sRHgh5i5LqpKkiNpG7uV0FT99b27ODXy
gda5BLwYA7+sq7JpMy3SdxnxjdBHYvSYpjneSZBSchmBI+K82372ZmoJ1jhFaQfWFGlPiFpq8A8V
dunkA/ijDB6M8dPoYMGguDTZwVh0o8jtlg3MiSFdLbuHbLVygtrY2vpUjUGmgXsC6aqmk/9ePBc4
ANH1M3FQZQe8Nu7eFLJ0sb3G1RNoeSRP6n3HiN1yk/o5WYmVeGFzdmjdt9mWqVsVrvK1BItDu7XZ
sRoAxEpPasbcEJCHA4hzSZeakVS+56mzvo3+oCAEvpKU96nE/b1NaWvRNmVsUVeFowIX7QFcm2Qy
2iEaW4nvSDN5kmskBxoDG8kml3TPtz5XX3rckm1tANUKj2i3l+RNG75zmSVIV4yAUY49MXIOvp4U
CngF0Z3N6cit06L+g1yV41CUWvy5xevGCJ4bW4mAOHmN2pcBB5wBDZ5oQRSuM5FAYkrUQvNvTAYh
WdUFkTg7eqwj3nNBsa+aCnMspTTvmFoTyr3vg1Y+I55STFKb8iDS+/bPmf78JHZbRMX45XxgCvfI
EayNiRX27iLJiCbWqSWggJijt7UYNPKKJzzCEZ+t9U7elU/19G1PrW2aqKBvQVF/01CCPvruBaqU
Ms/579e/A/ksB3vriXkf0zRGIi+BdgQPvE8FBnkvt8MFp/0DBynrXyvWgeKFp7Mhal5e+9F1vc85
o7dCT8/S2GHQygvLp64xIo0Px2VpYB1OnGVIacnIK9G/reK+8+YFV1JUKPljpb+1SY9UHvXtm4za
QeWb7M6ivMEHBDTcnOSic8WciJpfmdRhrjoQg/6oiNQUDcZIjv+COC37Gy3YQ+7yRAfd4pEWG3pD
yFsdyAL/T2ktWGw+T3Forfy77bE1g9bzCUTHLACQhIBwpFJR1I7sU0LHqriMt4qx39/vi10/Xq2T
lYWK2xAt7L72Dtys28TC0SX1Zp+T2wPIlLKOnr7Hj8fl+W/PWniSxWjx1Eck9jw7HHo60wx1R1Tf
Huv/LF2aZ8cFFQlE0BlvHQdG9SIfpEk8Cues9zlhj6McbZ3w1bLrQRePlPAr8awjzkAw8S/hz9tD
ydBGxz5DEw5IOx4SBM0jiyyuHfniPRu0ZrZBjL8LCEYNaKGMiSnq8nZkupVsvXevkidDt9KFWND4
HADVY70KL428CnDWfDG+iGkhsDq888eLqbUmsDUK5Fo8iC3hPS0WUYE6yV/e0Z+K13UHt+z5AVLb
3j07Pv9OyJC6QWo8lF3clVd9Xm9peR7+ttqAMO5P26QNsE60DZ9CLpgWSzxZfj0e78C9LWTy4lNC
JlWSM8q5zijxZzdCUHxOA0oo8CBvm1znr8WxB1tE8MjNyXr+yH36JkB/fojVe/+U+nvPVbScd0X/
r7pDE/pLndfk0TD1mckvjImJ/0rr5c+WS3qZjlZeVqozBLpDicZp7ZqOrXLGtUnIdOflrtvh2udV
56Z6qq7zQknWLwggb2YzG19amq9IemBpxKd26C8UH754VRwenElzwFcHXlI7wL+SwMKn4w+A5LJ1
4Z8EGXJ15isKuV69tj5HmPkcIXKeGVEPzEP9xRmo0Jgqfgv2PtrLgeyTvq0xwiy13RnQM97+r3du
6VCtdkTDdcXNjR3qChZg9nHOYJKRWAzSFZ+s+6pFcl3wLZiRQqWdU/gZjrSpLDdnK4Tc5ItW6NEL
25fCE/npNYj5ylYNu4m3gmemdDgZkf/Q9mh2H2OeqAtyAENH/o/M2l3bNg3Qd/Nq8jGyEhxUySlY
H8iMII37lg1RmgfPHaZUAfDaO+lsfcq7UWlAhmmIjPCJOIe+uRQW5xsFTFQIVVQgGaWRiQdYgH98
zzn6hi8JXVGZcBUlpVPscrmgcJuTpYUe1QlGTJ9+qubVdT02CSL4NBAq+ui/sAGTKKUYUw7cPpnO
cxktJcJ72ww2kvFkFdbjeR0AoSyXRK8N17wNrvQtL2tyZQrEoELFaTaHnTFmIeWwjx6wXNiTMxTO
HkSdcNI51/+pCPugvJua74hA+Pf5FMsnEAbAftcPMJKBfxoskRQIa37Q7RlUfwltVdFuuYndbp66
ibUhcMPtlER5w9rIbTYnJHbqUkHmojqZchAIzmuoWfaBPf1GnLShYUT3fjd/u5E3s9JOoCfOaSUC
7qeeQddjvMZPttl9g6zVG9DjIHH/Ximv+v9sYgVcPYzP7btEgTT5htu6nrjs3zuwpdtiYtZ3XIr/
MGT9DAZmw7oSbfyJdLu8Jf1eEdAOMO1JcLLJiXlXEEwayKyDIBk0jM/zOuLFMJkHeUqqjxi7EqzB
vs4PHHWTA6lM8Rp0DPK1rYDXXOgjVHI9twFLpsh7KDAvvX6eF8dn0lGjUEMHn37OfadACcWcXcnI
Jim/kpP4g5fJ9hCyfGAYsiUbhRkt78I3q/wonrGEVj7b9f6Mkb3nx3ZJAU2EL9Cm6h5ByLAFBJ/x
gN6x/tnIsOXQPk3kPnpogI1QGolHqs5WpfLtYB22m3Ta1DlrCHbMdL1iTTGUQkpsE6ZT9XE08hqh
g3Px1vt5XOk9Nkqt3m1FK+1woWVPV+GdqNtPBO31KX2fSOYyPPRWPviSV7ZNXrrWWpU2oikN9yx7
sVLqtA5ZcTzirb2OILInralkAc5gZ0wb07Segspy/EabTsx68r2vkT+1O85yIk+zoV/AV6+Re1pG
hKxmdD8S1EBP0tBSysGehRaxP9B3vsthNJytEwQPuuhkgSQGeVzLNR/6ftCyt2Iw45SaELPWVQlE
wLZFSzXhKLf7P++xmn1cHoVq3vD4HvAMxaxwvULs1dZ5WXkuc1SR5mCiPmOXZ69rnGt1zcyHAFOd
UmqLNWzC9vcAqbqwfjv8B77LoW01DSMU45yJnpG9ZF+9jNu57wCLB2N7UJ/ASTjyfJd4p1pBbv6Q
PhzCM5FbSCj2ME1lZd3TZkP3mLlYig9B4SXgRy2WDjk5HSiHnes6W/wdysEroGjANAh1oSVt24r0
482d1+PwsPDQpecil7jY3xSKmAJJJQ8pxGqeGwz4MjhuxWlzwii1Ia7u+ARtXjwhAFGNsx7dPG+Q
5OnPUQQRItIg1rRrvsmgs0bA8V39doCrluUI23rx8lKCOyOQ4GRItaH5XR5UwRNA9z3W2jCzoAoa
gQthGyfWjjihit20fVyskDbqN3V4Wcxf4uAI1WMD8S8Hv9CfpT2b1RB2HsVN/vwqka7i/G4EAsYo
FqCwDxjhiAkL189Ls0CJKl7+mtonec48BKlzqTRXFZSXiS4vbHEDF6RhHzZC/4wrAchZcLA4/CYq
NDDXzcMD+2h+vjyuPBNwQOvo2iZsj0Je/xP8NOA90iRZqw0P0oRnYUIku3nc+rpyUUb3tawBs5p8
o66zzztBWNsLWzezYPQXzVrClpR8MdJtYCJ9yG8aUyQaXW9wssUHPLmHtWdxdmDRleKsN4vgzp2N
ralrdwZSTiBGr3DtqNEOlHl67Xrl3NDvYr+PaccD/XIL0NMmXvR2q9l/Lk7NtFlsG2ps/TXrqL7K
KMuToxLfLLfGfoFyQ87kf99XyQ5ijZ7BU7ExG26ZQLrHVMdGbWveDz8fbbXTTA+xedhoBr/QvqEK
IMI7sET0VpZGU6TbTWNM8ZXq1FBEA+O0Wu6edWqcpn0xiBeBzfYxZiqUynQXAI4A0jRCI1CykkdV
QVQKWtOfPpNUq0Zrkxnu35BBPg5qzlP1yfAW8rTvHVRyDZWimYK3ss/0AydL6NEHHXuRGCVrsS+C
B3AW7Y8fZGD+nekFlq02Mm6ygyYtPGt6teleKcbNkgIAXMPs5PqxUgNyDBKELL/4iB1mrTVD/ekQ
laUDMHs2UjdLbXA3zeDxRtJWTu7J5fLrHZg3LvwGPCzMaqmH3tHcCbHLQMG30M+5iGPGkr0Yrf5V
rd1DKJWN0VzurOoMDqkFw734+dJhKgsn7j4KYTvRHKa1KyGIuEY6RHzOrSt9MEpGNAz3Dp8O1KIL
9+dIVelOktvJ/RPDxXHWn01EERgN3KmtzHM2B/6wbXDFaautIhy0FEcgCvZf6sajHETIgIRdCqfH
0+CyHHfQw79irSKEzuKbVUDO+6jMqlsenelrU7q3RAAGc07ylW6xJIHNbHJGoO6P245NhL3eU72W
kvL9BHMrDCn7I6AbtUMo78Juv6gwhREuWd+ZdgvwlPXDiH034es9DYGfrjFlovAUqo1yFDEz1B5K
Byk4XSiwpaGXkd9Z5Da1T6kbo7tRuxKlDEV1vbK/W1mtf1f8+rCtmG+8GH9BFAQlZbOuREWYUCd6
nENfThbJ3yj23oWS7GywLrpb8scqdGf4gCYGwj6cYjgYs2wtspH3HaY2ytKMdgddkExeGzVao4fc
mkX/wwpL9RRA06QQqSMAQnicF8xy3UuumxloIz1dh5rWA9LRuWtZe+7YipKZ2GaJD574zNmYyPcT
KOGelFX/v5R9J8QAQYAh22hLmQERXnad36nQeH+KNwA9RcOJtC/zpW6xg4YkFAmWRZEtbWKIrAP6
yo0voj2zRjXqZpTir2JT3hwtbJIccJZJLEDMIbni0iU7RHBVTEN9apPp93J84R3mlzb+HNXcrVQg
PwJvVVY+P9j6DXTdw0M81vv8tx9quQjCi/NcjxESU0truIGEEBLwWfDQ025bncd6uRAwkEh/+gse
4fWqW9DYQjm9Lw6urdUFLPVxDV1FrtgOkPzMSQETKNKJk2bBl9Xvxp5WgdNXv/ER8Xi8U9Fhlb2V
yZeBb7icrthYxSZIbyydbyRNVp8BUvFTYtg5ydlFPz033iIRQv2/twLW/z5gx7TxKR4fGAipppIQ
OaWUo6JGY0EN3qk402LpuT42VHRRUwOUJnanxtTgXiJ/DXLTz6JPHbqZY7AUrL/NvMABb2IhaXWE
0TVmX+8DrUGxtWUQp0c9q2HuKCz6SGdnFsx91hEULYKOx/bU4h8N9KuwNyWfEo3Xl9AH7y+nIME8
3D9OOU/JF0B1D137glwr2mQ90p4K+4oOV6X55f+YY7wak9Pb19n7a1rzbOxCeg287crLKFZ0pMep
9DxuF0Tg/CCiXR7tH1SxHBR+0WY/KvhOoEZHszWzb86/zfayORgfOE8XJGJINHpQ4l+tpPX3zakS
ldoh+6NT3QAdHddoU7t4ANHX6fQwTUbgALRQZJwcfVR23wv1msLhAeLw2gCafQtU3OSrOqcTIkRA
pg4nnt+NLCSxaZerMU12LBx2C9f8zpCD0gC/L+o5BO+uRSMbjKAfruITnuXBNF+aIYM5tEYxTQcZ
uHl73KUlM2UJeBhqCHSvPYtGiOL3wdS3+qCshsyV+9a3M0hYuHZGtEHHmZfFJ7pa/jc0/N4K06DQ
G29Ws3lFhHzU0ybhMeAMI7yAFXx8DUGHw1bJg0aLCQUc7/uNxYS/YfNLZMStcrB7+cp6ZLWVCPWZ
RKqBMydfnNSc24Boa8+g6HCagmXGTqnEwj9txgweez4hQi6oXu6IZFlXowXT9LiPFfVX9y4EphRg
9Ms0Dm+FrvUV/kYIRWI7OlsJj9NwyuNJ3m2X8E9as1KyFok4kPUCZrnKL7L7XIMsqxyfbiexT3be
87hyB73tzY3fVMU/UrSQq/rMsnon0N3rmzyVXlse7M8xgGmnO2Z/+3hefYUH1SX+FPlbvbmSNNdA
mWUUPxMue0BcLTIAbWbfI2qE3ZPBoMbCbiZQ+O/o4pQcGHnBOfPlkPB14JgqfIDEZakdORSOn65O
jhTs05YxFFpgiWm9PAie7mpruEGfMS5ByVsq1ttr3uMWefgm91L7PFmGTAmRgP/lIckoKgKTFSWA
Aw1UKQwJJlgVBvm0euukxHZuZqXabtWIoLG4CfXmQ6SzSKaBQPt+uu9zQ6T4L0ahB+Hq00zt9UZa
fpoAVsJZJLOh39bU2hzybOSDwQcdp1iumPKH9WJKJdZne1FXmAMO/XobhMrN401LKYuzreQRW11G
DfT1AoJk/7pbM8/yG5Hjdn9W6OsAOVZpuNt6CCOTuKL1Aeq2cTEBDSA+LxlqgaK0+LkO5mYOYiff
qPBqAuqGN1L392uaoPwvUD6xpywuvrMFUtD0gTKzHnwN7kIHUfqre9YkqcBeYZ4Lr2ecz9ucWRMe
cqaL1BARE1fOSkiTa3G0dsEqNLZ5v+RKdpu+mb//wpAaiR9vb6Y4pvwV8CA+Xni4rFddlrNtTdwg
7NXu8SBNj49m/JcYqdykkjGJqKHG63vc9HQKLGJvfLoBKMY2xdOHeMZ7xDdnBXxqhxq/H43EVHzD
R4Q0rUOEMC2gcBAAWAq7wha2SCfEbeMOznX7mx1q5VhNVDJUcOZJWirELO3RvoyXaaz/dj1HK6Jm
xcxH/BhJx9DGMFnX7hGNh9MvF7MJkV5F/2hW3vc7Ra7Csxz/fiKQMf6XUlQp3Y4eiMZzi8EuvoW1
2+Sk/cR9Mp9gKEIvdaYguCS0/Aecv4IS5fTFs92+kspwTsgSfepJVr/+edV3AlQP2pvxKgrtR5us
2m39IO7iQoupVKqVy0e1qm9kNAzAXmyk4bUh1cctrTPEdZoYZqy2f8WGhFjcHdAhLA0FrUXFoSt/
Vgq2t3eWG504LjsHqFTzLq0IDHgJ9PTc3ADAO04fCM3qkau/3618myr6uGnG0FXtMEO7pAqEBkpn
Fmiud6geeVmvohY8LO8o8rvkN1WVyL2S66ORCnNS10fqJ8atM7FFKREZsCk20/Ffw5NsRY88A81Q
/Rt8Zuu331drrWGFDkVvL7hn1Surh9yn/pjn5aCeOkqOatqU2IEYLz3k+C38ltnwUdOWgswrPsTd
wuRKKv8J7BJx3a0sEUz1AWEydR9MRMzyqzMGE90Bzj1yugwOHaTdz2wnaRxSQHYhKTFg56LUdvxQ
3jUlO6cj89AurGR7akicS3TXZjX3jym2ddh9tL8nF6ptGQIE0B0TIzyiLOKR2Yx/xBKeZPt7MPfi
vJXF4+rW0YMpDfsK6pZQ4Re20oKo+P6nZlqzChqlOHB3WX1lxRzQSUHEYdXHjPO0ny7exTwLw8m5
0IAJFnPfm5E8hnRlL1Z2CONaz/FBgx2+VCLcZ88ka6CEwiK6sPyD0SU1jHrkSVgfY0Nd1c1il1J6
0JdaezIgoZbUl5KJeUhU7lY/x8QocKWeUvmFeJzSVwwa8dUjEGi5g5b2QEnvDVMH9hHABfy7cJi7
WuKEXHrCpwVePWKaIZZhNrZTJArpUtJB1jvN9N7yq1a05vvWf7lZuPuk+DstAHSM01YS0HauwFlC
grwjiXEL17VSDRefuyUvdjX5xXkjqZJ4tu7+s+wxLzkPUiqPQalxusCFJOysstHaeQ1m9DvD0y+8
f0pl4F67ojeQL7vs+oVlfLliwwQ2jX4GWN0/WE4PGT9ewYoJ2RfoJosKOz2ckBE4hQh7avIlinOD
6zpoof0jVMXYiAnCcLs+RPVjABsMxdVVWeAn1t2t17HH+VCzVJd6iq6GYLsb/jHzbw0VUO8+qoTZ
sxNxb4bFihq2jyQVkQQEcyyMtFboH6sVb6gax0s4JfeVNDW4nyUWDS1y58jfQLrspA3DreLGAcby
JqEZjTCn5dzm7ghH3FcIIlj97Wo3qgOZnShYlsB8nrUtnSoHUo+fHpJqFQKz7C21zAzqxN6flHRX
G15k+qn0nuH5I/Am+FDCh4qtsuEvPTWO5AhfGclAZW1Onq14Pr4PoQjdzq95rZV1a1t+BIuZ/hwz
wIyMEWNq1+8GYyt+z5rw1zm8gg10QnSDJCuhqN1HVoafTBxwt1yhEvf+iXOiV2xBXYB2BIzhfp0t
zSH/PyocQiN9/7iMBBP3qD04aKD6LGhG4e99eeIOi7iFMqur0WaHswnndURNTJSEM0kbRlsmr1lu
3HbDy1uxO6qjyUqqQ4pqDRFm6c8k1ZSzkzKbvmi307rzvV0lUNZOZZlBisrzngIqwjxkn237tAUx
u5Nh1v58UtPJ1FBzrYCQAxLqxbYjsJLh1+SFrnRu4FfhshYQWgyu5sv7fhY0ErLU3HUQL/MPGKVC
It6QyOPyolFU3wQv3FPzKd5jCX1lwu6QERlg52hJUBvJuEwsUrg8WzOKNg+C8ag5Jeo2muTzIPnj
2ibCO2eUdWqm1xiLGOTH/In0agkYwLhNmk57Hkq83ZxHIgfE2unVymm9+B/CM4cTtQ0lhYGB6U/q
NFpAWGsg5/OaE+NPnhqJgYlCSOXkW5Dx8JrtwOesRNLkF+N7Z3pX81t+JqwcbE5EkzhQu3p58I0v
yaqhH4UtBcFgc/dUjpmYAU8mdlHqlddWzfxpKM+1HqczpPDzO17DfFolrx74GD9fYbQmO4CYcEl9
kdkhgo44nsqvR5O7+lumvgHPOhnNJvIc2aOdVk+1hopD6q6X5Ha3zQQrHTaFho/mqjPHuMbJzK2z
TG4iw3nG1Nkp9VLFJwr3G5U+jEhykxZEO1CvB2PexILF9KMqh6GK3/F9iUZILBYngx+g88KbmzL0
tp++cOszFgaV3RXcF5zBcE4QTl1rLu4qKcVhpRBitbKLuPyugToIFiSbrgv82XTfduCnMV+16fEr
10tPVEvGj3WLeIhKp31DbX+4YSvUJlwkr9gXdkBz/mDV1HXtzPvu8uGzVBP50XM6DWk+MLLbYXh3
Rs8hFetXHZRzQP/bad2J57Nkumvr1FMxoVa0I/O1p1g/MhBF1BiqVZotNhceih0fZHMEgUaDGfho
W5NPWyICAsYDtg8rpZtaIdT8FstJ84IqiWNqxfWXz8lWolZ+kj8GizqyyrhjrM0sY6j8ejm4syuU
cq3HvkyRxCeSY8aVKzxGOj4auk5RdRehUW+bCb5W0dpLb+5eZRc0e1/9r77EMHUKECKLnVUCFFND
DbYGiUbjP9wr+8tXaatU04F3K5uN3wgYW5+teb0MhCVCMIiKgIcCz8GGfacKjt9WuR64jEPxaICG
J2WKHPNdc2x7q8k1wBvzLS9mgHIU6IMciZAN9LxsThHEvcdA/KGC7DMWZAislxAdgEelrPQ4MTnr
uORQTIIhNWoRe/EvvaIImQgltzZ3vN3LSMSRLCWenxJqvQGent32hritsJGnRgVYHAAI8FfhEi7z
teI0NZ4XvmRHUSGidLKgxEHmcpZn7AoBmYg/GXGhjHs9Z/vhbSh0gd+6vi3xgEXRp9+N/Sx2UOLe
Lb3VGmezGg/OFnw+JKnm7e6zhGiVvZ7I07aV8KwYcmh7UmaY2Juyb6kzHEhbrtYEF0rC0JJ+FYm+
6+nkMan2A9FOTDAaMO6+vLb3NAmODZNZQdTFZcJp7QVmVWRn01plyeGLg44Krw1+yVO0BOvoobX3
19psCI99bMipAOAxZNpB8yegV9Ry7TEUDktpwUp1d7NKI5CGUWJMRQGwG+CITBI/vWL3tJcA4wUV
QUxfyXLagaGFY+KPmOZbOES2gBRRSdLz2uyQ462UOvtUe48nLSQhr5sQnPVmuoB0lYl5KT3M7z0o
juu2gQSfNhjvg03hOV/nv+78sHCnqJ1MYDvR4tnMXED3IHYOmFSXxetElRs5xWAjBtc1tnXUuI3m
OMBvdLFrkFE2IKGDxWreyKwoct9/iCIG1lsbdW1PIpFMMr8DAUqovGwtjOqbVAm8XOGuLTWfdZ1i
HWmpkN5OJRySITYdjc4L7p79heCnIwkw51WLyVciorwQ71EH6JqUetFKzIkDKtBiRnbjDoULoMlq
bbbGvK7WUmK9d9wFUrI4hkDT3XhxZTwgHwZh9/Gb+oI5+FWNFJ8LQyy9+847T/9JF63E1A+kqt8s
EljveJP0/jF9K1TkuM8Jywo7iupEtnzteSRpJ9qbsYDegJDb02vw7Qjg+QXNAYAk9phb0gZEZWRh
ZA40Ax2762lTQ+CzZtAV5BoVCp2Za218Y9W1k6rb0R62YubfgeJQCg69z5IRgjo3d49PTpV/7FRE
aKNZZcQFVm9xa6aLswP2VTOUzvpqfy7jpGmN0fooTQqtblkDqFUa7aWc6kYzY77Hlr7nW5iau5c9
bOtWHMvZry3Mi/rmzyck94eCiEQU0JW5phRQVmpoikQJ/OK5QJN6JMgSSEVXWQkikzBCTKFWfK2E
OND1MxDKkzJLNSW6sEfR+hdAQ2jiyPpYZcNnVl/4WuJoXJmXXr9AjoIuNfEW5B1WYfnxwT/q+okY
cf54giXA+y/hRQGy/vhsnZTciQiFxiQJRbxATGJS9q9Gzbl5y2976+Hy4bzLcae9xUhQYCYMwzy0
94zTceHYTNscdGBokf4AA2Ne23tCNdi0D7E54tMtYo7WilZG09mjlz+8YvqPi4UymzSC66W/9y6+
kghKCiObu7Xoura0Cb/tO7JmctuqFjAhqA2Cq3l8xwC2D35T3P3aD+Zw8VElFk13D1NuWiMlmviU
bZGDwdiHuoAvksQbJ7AE8CwiggvffHrKT7UimwZ/k27mItomXUmDSrfvTM2cWQ3+zEMH4plWVWuK
3HNapRaZdZ+VOpKBseW1raY6HqHzxfmLz1uyL2I6453PwC2lzSO226DB2uFbh1AyOBcSLWgVQrSt
m6Iz/XCRHkNFtpWVHGg65RqVQClUGuPtYkt7lxww5LtmPaDOVSGwia5sPZf+EnWAFXzysBR67USF
GSY5CcxqJUOdp4jpUaPJntP4d9Xw/5PYNCVx+P4c9qhMbykpmeFK3aF+4U/oIsKN5vUS+1//n1mA
JpsrvX2rlo7feUV2DZgeG3SRHbNPq4cRTUMW8T4NM2Fsadwchhx4KXuDw7bH+2LUUl/TEsYcCFCv
BprPez+5g87kpHTyetCaqpFa7iBngiBT0WsScowxT93GEgAVysP/oFdW9duDnccep+YU0WxAgrlL
W3533FQqdbbe4uG4pzf5Y+j8eUGiI4HAFPN4DPuRAklVTS0e22jANXNAQehl6ijIrT9/Y7NmQU21
Asg2W7j345uusDKqtVc0lXsKGjCVIcj0BNegswDZ47RtQvlRhiawXC0rdp7IbdDmtpjCrPMLwim6
ccxaIQypRgrMVOpuj9n59iDPoA9yQaffAbOYr8vupBrcR6XDvrbvgjpyGRUAJKktms7IofggEVXU
WUY17u1LUW2lwfb9XGtAROLgv0VGF4v33ubJ4nVNLtoWd495CwgtCzarxNEsQrgc7QNr748MeBbD
aJJ4H610g8mZOEdHbI5rvShb4BaqxqawoRfiut9xLHk1fKEUmroir+/wx9Ag3hT8qnASs7rzXeq7
jgoyWHat988cx9fXGJv84c48WeeM9RJlS+AaHz+NFkwug6ujZ7VQi7eV04Zyi++Jf7WcGx9c4PvX
j2giKmD4WgLyk13fUn9Q0z1GJX3Y9lH7d7AOaNhhKI9BvOZiK4C95gF4MJc/qOWYsuEI6j4fp7Vi
V6BHnWM1zJTckNFUKcGr13p0WluQhhRHdOqa9pmfuEVSfzwUATm1L94t3sHc1pFesh3fYQBDsVy5
7CpPkha7KSs+e1Kljh8IMBsrpczhoKhxxyCGt3tJaFFFuD04Ke5HmDSrTcSkRaI8cc++edDz5gfF
wW/wM/KOKMylS1ZnAhfFK4d+uCcZEUujU+42Lil4QVpkaxDJMv7HImaSjMuwP+g2UaoNyEqY7iIO
YRkQMqc/317tDh+15zC2GPAO5SOyyBBlObolgE6tu2CdV3ukI46PnNqd0RrUswcwju/oF3cwBtBW
rMjGICZvo1xCMt9B9dIZF1Ih9p2ex+z3d4EAoKBJIMeKwm9YDR6RukprLU86EiCblOAS0PlOF+fJ
KcGKsxH9dwHWkw0D+oyrp4Im+3SHcOzfF/ooWILS3aAb+UV+DcA9qMW4itDj4qH7tSFWpCR/9Cpu
HD6JRdiKg9MeEQQn+WhawLo1y/dDEJqMKEwsA0tLTn271V7Z0Z9ccxnLL8bqu2DU5i7Yz8gLsh3V
HZfOhpOoyd2abxzIQoEKMZ5M7qaMYFEPzORElZYZEI1LGuOMSYgRg388Xq7YC9HvF8GDlxish5WK
Xn74pWDxhJSu/t5OUQ9e0yNeCn9HhDjmuHtPtvFcImjiHGa6EVCM66bf0IbTBNbo2Mq28u0apmxh
AUpH1rbd/1tto6pkwrP3ad/8wiWkwO4rEYwgNjF54pnmhjqiDHAfzJUMkzdicNTTFV/G8lgVIHdE
JBw9hkvPxsUKKKo/XFZ1yd94XciwWc9VxUc52BFMyRdSfvTkXdeyoO5CTqUfDFFw/lQpR58dt9We
J9TmiZCkNmysfW3FN1yy4kzxPT4Sw5mKUxyjIK8kShQh4NMjjGIGoVfYhrw5bYQ37RM8ee5xpAKl
6Co38dn+qBU9ZSP81GtGsn1zUiwWvqCoQvpzYmC++RLEooVflg+WRloZX3oJibaZVUlluR9pqu5W
UpwNvtfwRLjk9cH6shK5ROC854PuRACENLj3/GvQF/cTiWl6//rACaUcbxM40yC7bWQTBd7KxNgA
WzPzOnRaEO+/beQ3ypjOD7K/Wb1GkYtRVQi/nT5dVTR7g6rEWcAUJtwyxXr0Y2xXqRW8wYCuEXhO
WIJ6uEeGJxY7uE3WeTcD0ytB1rvFL64ifMVFJF4JsdWNkeXxGlga8pWLQPlxZf86PUv6g0lrPJhK
LdybFGXrDOeztwUEzXYOvotsfvCSU1B2wlCp7s91rtjYDqeuoHtA0Lhznv0rtOzbnJvygCTWrJXc
tP0J2AVc2q/Pp82JoXbTVsgCQ7QElrYXs7tG31Tnx42+cf1fLV5SXyqLXfnD3vnxyORNHjSz10ea
W7pkk2Twid0Y3aMFplGQ7SzdXheHC7uyu9d2kJN1st6xnk7jxAzA3zJihHLWVLqwmOJ7wiBXsIkF
ZGkeYyk5PJl3AQin8y/P2/OmVnybl+17e68uLSZ1YK1tF1l6YGjvwW5orNEga+Ydqm7L+aj/FhXN
PVyd0C1173lAdgiQcvUSEKv3Jxy28d1O5SNnnsjvt66jtBGR+8CSzImwAEA9HlEZ2P4BTsKyjQAc
3vBgrLuJbENm9qqM/s/LLuUoewbkGAW95MOkJ3si4WNVqA+QE+ahRGFBX0l/Yy1uJm1uOsqM7GyQ
cmnVSX7lQgxSYlqf4JbcYsjHy9zDEWyDgpvsVFZzZhW9I0uDs7e6ngnIm86LReFujSlBQ72e/UiX
v1VtRzLsRTnj7iwNBUx/MD+yGOrgrVwgsD5GEP8DTOJ2U9V0DKzFuv8Cykt8/cJc7johobQHdEf2
UJk4+N4l1PmTpLlez8c0Kxf9XCvF47n4XBdJ8alfHZFwXeO6tFohw2xnZgn+1zahzz6hebXgjG77
9Zdh7x/3zkZX9bDb7kfJ+Q9YZ8RbJxPuI6QwpaR3vG4VmepbMBy+yhef5jBg53uKf0s1Lk5JR/e4
ap0Uj3capPuRlRZVCBzV+6M9887Hz0HIi+0DXJKvRsoxVuMYMwKCfjegeB3EeFYUdgwnagKSu0yx
+BXgHN5w3sFJh9+p6X5vbFhpXzUirLsRNMYk1jPUKpHdkCsL/dg0bnbsrwUE08J9p5BGQImwBse6
pRwMuQtxe0iRbWGFfyXCX8eNdSFg4gb7cXSp8KAdJAduU5MAdN+8FdYfslkRuAC2ePqofesi+2P9
94i54L+aR5ZMzPeK3tdXfOngEJ2thAtBNOyKJBVBs46e1xaPjeo+IvEzH29jHW7jKnIpftM08Pnc
dTxCx0LUvpIFYDKSoB3UhSsU8XLfUEtXU26fRXtRBhRt2Xm+pr5G19Yf1owbeWblyQ6RdywYElfH
4ih1LtKJ3yqCiclEkTEEVXKnPqHVVi6bzhDQLwmMw7tDxi7sMmpVaMyeLCWF+RXyX0QrN/Ss3GAI
4CFIwsH5F6XHWq5O4P4Cjao/htKdXOKgQ/DnkNwoPMagc76+jT47z+e5NzScv7HbQDw72U7IO6zM
DX47MgJrYfpqW9VjfqEXINxhM+0aNGFPjTgEXTubDW40OTlD0S6BjHoMOCQyLVw+X9MFNzJPEXOa
mjCkmx4Hs+Xk8oIPurcp3myAI/kL/wImJ8bdaDtEU2eZWUoCF+3j+5Z8FASgmPci5vdbnhIdVfWB
Px62S3ko9zknUQdz5qupb6mxBbqurDg1GlqpH9fIqChc9dbn4I6Sdsal3NSO9CtgPsoQPuvSlr3i
67qeyMFsEE4rrOZR0WcdqX+4KPAhnL1oGGhCUbFGIkY69wogLtezaj4bvojdb2P2/rvstB5Tt0C9
uigy52OlpBD/Wi8pVNM/UwTIMwqVWqQiNwaC0ENPfB88Eq5UtMlC0bny69oUq8XpQ9dk1keLWSoZ
liaJN2oYkd8WqHgF7upcUjESRNlbJy96bVb10oAZ4hImE9+Dcm20DyjhBwaExJIZBvgAAY1EErfH
sR8WR8xwTnYh9cp67j4zNYjmyo6K85pHe8su6RQpqpCY/dYL6X2E8eW17570c+SzkRdycknPFeP8
ucYTxW1vsbmi8Dqw7TLLXxvh2pp6SIMfTCyPj8+d2gS+nvjdXu2zXR+/xmdFurtR7fyUS+kU18T3
3QdzkpSJNl1bqmQ3XpVf/tMGwphuHoBl/jt9GdEBDqP4hk6nABS4YACE+umAthIBlZ7HUyBrtFZE
Q9ZM2x4HV0T7QTrhCzFiqcBCAunNtcSfQgoivB+VulAOvQ6s9ObXoHu6UkfSmjUdlPNhp9Z6ZooG
+cIOEqxMZXYdcbdDCqovhbSUrOtPPKYzehkuSsN4Vg6PxVyl0BYOSm0Agne0WvOZVzI6WVtRwk7m
pLu9IAIPyJ+x/FF0Dge+r7nF22VU9vHuBpb37tyjt805Sm0E0VOLIPalUtmAj9n+hSIpIeMLHFgk
JxAi+0qu91japmIyR00/24VcKSW5XCZv95R+kc627Wr7JDU6kYMbz0LA09yeNtA5Etwy73skzWFf
JYUnXEH69Txpzci05cvkqadGdwjXuHyi78bVIjzTxOfIkh0Qn5jucSWxo2hc/+T4am+KfB68idGf
l9w9Baiytxk4PgqSAeksOM5RSsbBcn1T1KEhQXMJUXhiM7xPlflZjFthKj0xrC8jZmU+BHkZwrHV
zBgnB5GGmtx0baEYvqaZbDe0DxE839XUPdG95pZXLxQXYhugJsIliBSfetG5jM6VnIyc5ONbnOSm
tIuvxHwrSXtSbfM0vg/cJJNKisHiaGO/epgjyhHDwxR7SrJYSAsRuJk8x+DIJkETU2IxA6/0JNN9
68G//rniz3aY/shJf01BetnNfB8jVPpOhWTBC8LM2BxCOqK+xqk+zRBGz6tlYJXOsZRr0tx3MII0
7h7a6oHybscIRoDeJZWISNrN5kK/0lw5wisnKBgmIYl0eFPbi0Mto65EY7SKcw98vdO5R4AylvX/
sZKIbpLo3w0041026j5pWi41WqYwjVeoApfaqjSx4WuCYJ8/vBO0H+1l7496G2JjywcQCkWz2OUz
ZlyHAmA0F8cugYzVLZ1C5avet1ILEzC+Kc/mziZH5pfcTGs0iE2E7WxsRtEevcFCAdQ4SkigpL97
nJm6S1yLiajPDzL15aupWrHIIWg8WFYgFI4X32wdwkZQOJ3otlNYlc7CMIaRzpXp3IKPXPVATfMe
VSzS9iEBI4aYmG2Kw7F9EtJf7+CtOE2JgPebRvIbow2QTdKrb+5ULFRfTNV4vk0nuM2toC5jBW8W
bMDKGun1XnyHacNRfkEljmEoU5bngv6sCXk/EFBVHehsv95x8bd2P0yhD9sMyGrsdeymnlbrSTzO
n2i6+wrsNhljJPky8nVYXd9gk6ufVFkeBVZPCq4sc8fZQhGVO8NHrhBMSGkdrj0sz2XlS957Orwz
V3MTB0zrFtJgnOsVSD3KD/1Obj8g2HYxLPi6X8Rj3dqKxacbAnrcghvgFxqAZvu3f+R9lOMa6fmE
QBuJ0WEwKBwVWeJCAnQqzJzYWJl1WBLyjfdDlt9/iyYtC/R74eawRpz71KwYvepeI+VmXVq1BXQm
DH9LGGOLpb6DXb53qCvwkXFGhmcLPzqlTa/5oQIZxYSJZ6qhFAyqkmXTKUO9eD4tsjOS/7I8LQ0m
LKN23YJqyxp4GozSJsd8lbJ9yOhLWRMlPaBdKfHkyx6dA26iLd8HDyYl1oMagdwoQyOPwQMX3h4N
/0En2BVAGkdcszDA42RstwwoOqHxX5yu6moNhDoxTSNDG0FDi+5GZRZ3zGeRr2Ta82Or02utDgsQ
pLVeQAQouEUlDhfch2Ks31Lfv8MIBT6FdmBNnbAjFEGLumz8TtyTFADzWS9pHD1Tm0b3vavC0zgP
0lt5N8K4B9efZFNj8X18maoyUgfTnW9RVLWWn60TDUcoW6fwqBtevOP4uLNu92TiWLQ+dYAsFXdr
ATb4f3r9fQzy0XE2WqApzbMZw5x9XSMQGcWA9XNQ1YY21WH6V2rMaTSbVzpqyLehaXF/+yQ2PiPW
w7z+gWsumLtc6RobG30Ol4MNnuL2/+fGi28SL9ohv46gIVry2VLuRvyL98/xHXU10xFNp+Gp2RMw
Ni5e4qLefrBQL4rGVHMpOX9MGAsgBByMQs4HOsuNj9HRUDbi1KmiQnAPBCaX8LsIVRtZsZ3+s48e
wQy+TZ6y+3E4DV6ckY0frIJNt8z9X/6pztGwfl6hIpnN34iKu8mTpKFRp8UmWrLs8UQoDVhcDY+N
vGeqV2l46AMJhQC4cTBsaE7Vv95UJBgnpJjfaFVqCidQVWQYAf0W01GPkGHZI08i6vKa+Zx5eSEW
BwahbshYTB8BsUBHOvgXycyGBecsdQEKVWjmzknBtkrvU1gKXH10OaI3OLd6NK/z+1g7xaSokByC
2byquflOmtyeA6PVMfKKKGZEYLKi7hrJv3hbE6QW+OXQWNh8GPc2uuV3CHAfN/XznqnC6r4z+Ex9
ao0j+d4B3X4ZugRMRm5sUG/Gd73bW0pZCAouGBOZ+wVcw3E4ERt/dkqbmEaxLErbDAZrJUjvHM1j
1e7vN0fhuideQ38ZuTMGkGO5IPQffnuYVEOi5a0nEYr0x54jc6aep7oaHzp3EFu7cAxOJxr9EY5o
VcNjA7imX7w5qj4E1z7OUPLwY1Nv/yqgY2InlPng5IYm6afRfur1J1k27mdqCzLVdclJNbp+67jg
NX9qh3SsL4Q8nyPgQpj3bQES0aM9atAhUR9g1vhiWIkYlxSK21O1kqC4llWDzB18UKPEHCkOpVlX
3k6j8X+2gys5px0FqGcbQHRmgomstdJ2HlqywXKiMIb/CDmSaNnLVz72bGtTlxl6xbzTovwM85dx
iYgaVHHk4aj/tqDecuw69RXQWYOUpaZXv6SU1yK5FTfmS2UbGfS8syd053ww/dJU8PMA6JbUbdD6
Qyl9AidDJJyQNROic4Fod3c77w1Bph1HdFldG40KFhlnO/W/Bce8lU+PGyD4dwnec8j4CTcLDeJv
ZMONgaCTskkx2kwovAMFR/w/4NPgVVSSQGh8LTmjcHdZsBm0rxwuQyl8v0BrdxY2d/Acol3miSip
vL8E3bq1iwx/pJrob2ehEMgibzFAgw2+759zdMWSaYgT+UUk38ffrE9btt2vznJKvsREI39RQcB6
MaC/jXfo4gpt09Dp8png9q9NeQZ2bpb/nUHXfWPFH6PizDPOr+OSLMFr7fTDGHATAsi/yP1yM+zS
ikwzs7dkiEgqdnU8FW9AGUtDYDpGXRJ2K1IKrSxp7dU0arPBx6mKdft1XQtOu4ysWQoo0XD91Y1P
Jweo16M94fI3NKXMXHJEu+N7NJU+v7YOkkkmyEJ/FAamT2cRZEUT11XT/xvXFHb1YOds8fXf8Je2
cJpve9cvaGeV2/uwNr2diDL8eZDYa970lBXltPOTAXmxkPc2hZx/lfW7KMGesX5miYhjI3UQEptR
UQbQji9VSmjpHxmxmdvokp45UV5bRSZI/1Y7tVJ0I+h9MgJQ5codxV5y9o+OOzImlc5JTVmbyd8y
1aEi76nZvhGVLWiS2Y5BeFIeGwj5S9sexCAeGTufjKT9rQlluoEsK0nPG6ObvZ/acGDUFpyOdTir
4KuwOh9KjQUiAAxg/e5cTHohWQ38xB8k6/jrANhY5IQbyVj4Y8CsHevF2mnktihc5E1L0lrUkJbE
TgsYK8P4wUbLSo/RbUkDd2pjEXKkN9+BjQx20QMGfa1gkkEI1VbOCy5hZagUqnr8atVQsGsm9rRE
ftuM+LYoC88OJghhfRj3PeDniMbHG6Qxr7nLdpGlGgLweM23BpeiF7ewJMBy0r+MKq8IGI0YSBh6
Z/i/Ooq8joFr2fSTX4H4nn3Lz51i7fYUQmqn6sYPTY5qRKwMrpjNLRD5HDZUXCGwa8z4yZrcZIje
OM4T5VbTte2YXURljIuagGMqBZBRnNW94YZVadS7S5TtkngFaUSAlZJNCnHLiXdy3ovH71r0ombh
mVx3C8xfCZdfHcdTE7ANx4kdh/mcjkqV3hKiHCtxFMgtXsc1uCCdkxA+59n/nZA/rrTdlWtVlvgc
xOJWVTa3EgrYtghAD+1NYbjxEzgytO/43Owi/5lpSD2Yd4EqMqvn2X9LUzbBvk4JL34AciojYTCO
l/5EZiAmArz0bBU60tAC0iwWRfdyKIOs1cNcDUaP9DB/dGmktfvG0igM1kIMYjAMu5hne8A1Shvp
PQ9wQPgZEfkaE4TwfyonQqudhjzCDFm6vDD1XRtRw11OGlA0akimEBoZX0gmcN5nDT8rJlhHGHwN
QT8YGQ/A9WRbxd0Xh4jEzL2bYQj1Ly09H4SBITge2hTwOwso0iOaX/ywhg4OMTezMBoGs+Z7yEah
fTzCcwbOvVnOPQyOEz7piJkZva7MpTR3FNRpr86kCYQF/zbuuswpnDBSCpfVBU9fQHe5a68goW5D
rKlySpKc5MTvE0eo4MT3oP65QZGoEKDy8ooaKsVi3/0hbqc4XadeHkBhCq1mXHomTsi2x3D5n549
BSKfW5wsTBU0sMhLfKd1WmBzuTK7yIdH4cyqpYVFdlpHphT0jzZNwhSfuNbUv1OzXCV4y9wQyoQU
InlM0phlhNOCO/Z3RvXDO0X54WlGvxl5MOTJwqHE+GLybPh2hMG2xG5v50HxBIPuhNk1fzYVTm2D
FcVn2TkJrLlNUuw0FMPVQQIsiqmUwxidTzOx4fI9EtW96F9DvupiJ7Mshxa/0AgfxDkNL+nNa5Zd
DTPIjXFfpKb+PxVBKGOW9QPAMytvxwaR34/VTKEoUkGumHHlEC6RIII0QWkdXsRYWW3aJclg11PK
KLIGWqJ0tsAPnEAC8WXjuqFl3pAlS3nj/u1rpLH7eeG7RjdvERg2+byOMV6rvz9yHKvfRlhd+F9M
RulnSq9eFBofrcT35BKrrVUrxyZ/3wIin4VJfNffAsoEo3mg1ziYKtK4n48xzyp3P3Gpif4IUOHk
dV/TNBsHoEboObTkvsVw0adM4+Bhqz1Rn8iC1fGfYMjJyudgf4Gt3k8b931U6qM5Hlp5t5Y8kM6w
w37fKJq30bp8vsiD4ruBd39M0r+/WiCq53YHrr/duWuWa6iiOx0Q3R2jb4NNpSi/C3NJvTU6v+ir
BublSaTBx8I8ak7K1b1po7ZG4+SnJycme4tPFLVHRpBade4Wwqxl4wGUDx3vXhUIvIJcY+zCg18K
o1ghZilba7OnebEJlFBWKKHF+iWLLLfyZAxh2yCfp36VqowbgRcn1AHRNLlVJdR5XEmUlf3M6MJR
kuSMmA/85Us8NgKUDC9IC8ACbYngqzVnPXo9pTXC6uvdnhWvukE2T2CKzmySdJ4XOvwnymaI70d2
e1HtnbB8TVKFLDgD4oyp6u6OSApdT4UQyj6f71I+abd2hIOg/bO8kPW0Z1laMkXMEc48U1RHspIF
PPsfYT/PPV0JPksxMeSUkMsDeoRBTFZXOcvwM+5lrDB9I17423kus9XyK+0q9ISGWrybafdOWFPD
OELqheVGkWaiidLNiOy94ShPlcP11MNO1URgRPkWvmv4t/a6eCQ3B1f2tSxBu9wHiTZX3hCUKv+6
pLv7AsLDwhl6aaXe/boKTiXB5qqhyJGoavBzasYz1rvY7IRBNpl5Rl9uwBAsiUzEMeA8Jx9BK9PM
fmPz+Vf0l24GHoo76flvRJ2Xxi+7qKG3Bhhm9n4KXpBI69Tzxs3EG9h8hR/dFSJ5/8PEMS3kE+1G
ExS/zFIwYy+8tNbA6POrtgzKe+dtihWiQGJpqDgbEzs0/kEEDIryearEJ4m2PtdA9mS/dNQd/eE2
IZiyH8pz9akl3ZcBfMbFHngSom0hj789Ez26s+aB7MSkMnCEqeZsWgx0Uepq3G3OOooQPx4kvimE
DuAXLsBl8DfD5XRHq79M77gdiI+/9DlV+fD727xHNvbujsI6gfgi9XYnE57OiJPd2AA67BnUZOnw
KaPu7vV0rAP9hQggNCVoJHowOqMpYY+ew28udCkiTqQ6MswIkxZDXPqGu+BOGjLSot8CbHE4NuED
3X3rNaPfdBpR+9QpQ51GVIwOe4w+VhgbBm3lDzU4Xaab9269NdUeSmMGNaBpXTYv8Ok8gQGCTbuM
3NpnG+w0P6sekzqbCjYz+vYeqVljrFwL0HmEm/au2N1H6iepijR6H6PJnmCEw709+rgVOmHzlnzt
MQ1sQsQIvkviJwC6csoaGtFoBY7iZaprHfLXPjitY8L7qwEcHdCE8NFom1Lbs+8/YI78u0rt6B7l
qS6yb6jbga3E1v1YRB67GjTTZ3oEvAUlkkrpjO3hJQcbEeZBsetrENv35+DMO1FeQOtfLHZFiqv6
5krGzbOxwJKp569gkBUO80jhvtlPlmtiqFxVfP4Sf4m4OltXYzZjYte3XE9wephH0YF97N+kP24y
TpU0XxmX/un/6TWetlbdVlWZGLHtKco46yLCmSi9kr1pcJpu7lclPVZEytuYlfDbd+rctXdt6WVr
Nq3YadGPGn5VtUQ/gREYRF28zeFJlOYwsK3rpdLzZpXMUR8u0Ip0TvQcX9DzcPar1I6AjvQ3vqOx
6VkkEfHw2Cv+WR2AZydplqduWAD/Aisstl2EoMtr6dINxYSJjhihv2MVAtBhvaYbHCwZtlrTFv8a
NnralqFCV15mxWDy3IoGINC1KsD056UijrDuKP8C1vEachppWW3Q5z+1xHJx1Q/V+I/PyD5w3+9B
PHTEpjm6VqrZZku6A+eh49J7VZWiE4Q6ebMhA0DJDkcwmpCRGiSoqxdpy1qqUJYzP3oX309mmW2i
LFwHn5ngH5hwXhJtas8vjK0R070zwAWclesQwkEHN8h8y0fpfnL/Hue3x6/WWew4koV6pL8wWSwb
pZunhlf3pK7A94Rj4vnd04yEkaSMGVxeGPBuiD+wOIrTI8nlZ4aWkvnKXfHzQ+OK66+61Sv4unSH
IEy9RYEA2nZOEFS2d+o2faRTTwPun5tXMofGzJR+DunevMiiWHVf5J6F+eRwLSqujZUO72Yt/KEj
qeLPCugKPBjnit3Cs+os/EkTLOOvtUkcffmdYeLauGNKlQVfk4pL4lnK9HZl7tzbfzoXPmS72WnA
QYQkz57y4WJQiO0G8q7Gq0nIjx2GclEuReegkdlW+b2pDbbU8xDU2sMS3wScm5O8W3oNH/RDZ+J5
DSNOcpDAUFtpxhUyfq+746F+CmAneq+RPJHgKJFoBLWzMsJKYJT/eNg41qw5LgJrywh+yCg8VUgS
ZGq1WorVhU5Lrz2c3AfEQfzAPP/JCU85/9ENK94CPqGhbwSxQS9C7cKhuMxD4l+ELY2eQR/AbCzU
VoqpQd6ieqnPS1I3CgnamH8IWmG+uG8/9qUMrFE2SPm+VLh/TzKEee836ADkVuRtBMenM7JAPIL2
LeGxTw54pWjfdWoinNgdLs/vJNcY5VoSZOJJmTsXCZgpD/LbNN3dTJ/l9oaiH7YlEdOzlFd77+BA
gKOOv4cMawqByVxIyE7dB4iK4y1NHl3puqezG3IWVTzbOitVjfLOpfGw8qvb7epRnnjjoF/7dInH
Au4n/02uz9XqUxVbDI3pGi3Z84cKPA1t0Y79rkY3baKRPSmU9NtSddLH4e3uv09zkudC6Jlvx9jk
ZV4c025wrw/xyoBTTHG+3Oa2SSm5QDJfSKaHha/Yt3c2WDCr4RbnCiSWWFZrZ2/qCGXIx8LxZwcV
NOul1InQjyTDgb0hPAYiAW6md61jOrR+t9AqyaxSrpZ0PR4HbV9Kbxa33xmvi4z1xD+HD+VgfMEa
2leFcN+wb00jkt4JPtJLeXJ8ysLXE031wQMvWANqgEahC+IuN2Afs2KsVWDLCWVgQthGPz6jmvnd
9/3w+ygY4Tpg7SQ9k1+L599HL0MWbXjT65Mehy5w303Koe8qtG7DpPKZBvoh5MNtxKBQugOHpfgZ
/5M4GUV/feZen2M/OFgmMYtjuSQctxOQnqjPdY/PX6v4YnTWNigG5RQTN3r1yVO6miybugLeAsLA
TFugSUzKXU+Uuu5ovHAE7gaho56aTA7IYtAnTogH2zOsSVrtiCKG8OAGoIIMEjKPUJ2xsiSu+cg6
ZNzbo9E6qSW0485uyZFyuI7+lsPFd5fmpEK5FpwuG8QJRZN7RfjfrLPolXnnAjgVGk0mxF2Zj6Nz
pbayOWJCVmb3YIwiJObvrOpJMvnVAdFPgrI3A400KnIEb5bAHHwZgTEta2F/tTAl3GNbV8K8gX2J
3+t0kfiNuGUY36ofXN+T9s7e9eV7I/eOOqJg1gL83ixGSjHcVS+OUuWxjRhGArVwgsSk1YRXKdbW
S+xS8L8m3G2eei7XrB042MyY1uMdNYBio5t1uYDBmWwVVUbXadRz2dLQaAUATNJWfWu2w+J65+5I
e7j6aEbCZtWOt9rChW64ihGPopYzzonzF554leaVmCw0JjUptbKS1SnSYgixoNAJqIMAe8AswQMv
LXAFGsEmrSU3nWhQ1gaeTnYFrrMos9RF5b6AzQgu/nMgVv2xPDcSzFTv/+FfHq1Yv7MljV2auDa9
S+ZACv2KwRZUyWMCiOatNlfVDcXnZMbDSxwKH+NMSw5Odx3Tp+zk79Moi2Ns7hB1wuNWLl6v/0f2
FkYAFFBy39dZSrNgVDXo55s7bwQYExlX/0etEjkQECR49akj5uozlXMyLNHArbn9T3hmquRCbgjj
6TimvLnDIqHhNWUQFXQBAuKer2JP3L1V7FoAkOfnijXL7YvGvXUzyzqn9Pbuvcp1EmrYnffFngx0
zPs3GHtomBclb5PrxI4K2TPg09MsJubxQSMiChC+eV+QNa25+sfOWk1Dmv1EHSpweQCvt+yF2S0b
EQekdEiiS8tjG5o8h6aIcwkh1q2yXk9Mf6dU+ivsnSALqBLj0P07/+pQrMHts16TgYvCCpSIR0dA
1m2oTHy3z+kPJ6WUer/4hojk+5534ppN/sV96D9yyV/H1LaGj/U6s8sWtHncyUxwL7um6DXoTKlR
LBsgdKj6X7eWo8Oy2F/K37C6CCJ5q3ouxq9gkRt5uuom2KSYlidy2CokazzTOqG8zyLc7ZnKrc0B
q6QXqPW24sx/uzrmfBbivalkwSIxGI//vkoB9B4G287dRlqf2lmT+w6lxBNPHzU/HOE743xl5j75
ajRNdd1RdP61ZG8qmbomAq8N4sWolNI4BQWP2Fs5pcZ7G1pk5zRCNSjoxogPnUE5lcyDOOD51Djw
FkNk2xLEYmaYCqpOhwivtv8CZyO3CDsjnGz+YgAuMeD/GmDmMIEPfk0dfzU/I0czZNIk6L7UBAYK
KgHmmVv0HZJdXdR+3l3SofqGS1rIhLydGOtiPqhxBbzWzaViTgl3g7H/X6N3F4/gsUC8HIBwQ00W
11RkpklN6CHPCID8ukMMC8bYbDs4JAMWHqLQT/YNk9sGY5qOhG/VOuopdNa3pJK3IbtMeHyB7OJS
P2QOrr95idpx20HXQunBF+OTH1QzEX1Oz1+Ha6+9ZjFzqclYfQ2HXY1iowNMKlatQeK9l8B8knPI
rha/8UI220ic1DCvEDp8iEErlFsxyoeo4+zzWz7E6MDoi4tOAuu7V6aLpp9M2LgVLjlq4RXBfyvd
Zu/T4YHZXDq13LdTcn0BsJm5azImn6tX6mtdit+4X/3B1JhxXC+RPzsfMclpB/iaj+Mmf0NLW3Xm
UBLKBHgo8/JCMgLPWzP/bz6jSqOJ99DSXaLeEbJjPifp6WiwZbT/+MloOYKHuVgU73z3kp+bnDky
y93zqFKzXIE7wIeyphLuH0ecz/hdxz927sDY+UDG0D/BAN211KUYudoJr7TNm33POXWw4oKDqqjW
UVwFh6iWyzB1r+G6HtP/3r44oxipE3TSPlXJUdKuOcFDfPCxtqTBm2VU/rvAfQB8J5rT38J4xyB9
MgpcVRcnPRi6Y0pJ9+LrcEbgIm1uDKNwnZe8RJa1+vSE9L7dzP05d+p0Zmu0UBRAx9Ijz1O7sCC1
WFViuPsFBtqDd3P1G5CJr0j1xYGsigUqFYXnojrsjfUoY9xCG7hIPJa47zUScq3zENgqCHVztrHh
t66JwZCd9Wb6ICa+YdXIikfk9BqNDtXswL0seWKZlj7jwPW+/qlZ9n1AH/vszgvIgBStXz8WAUWB
9J3dICCoWZ9wViaSUoX9eQqMPwMxvQI33+B6UQMPOVWx6Pq0KTW5xHrO60ESMIkbL1zwfdQP5BJD
FlI2Vx+hlOA6BofRQ6eMtVFaulsfr92TDLfuNg31HbErBrMQPrswCurmW0+rVrzth4GXhNqQhyOk
EVRv1IDzP9IrYG6UNMoD43RvZ8y1eknsXKNa6NXmryu83DPo/r5plMBpOTFyyi2FW794P3Z9WZfm
h79N6oSgsXohAHoeA971vxU6BHh9gPAkerWzben/WnkPkkX3aa+KyUvcMubO3G3pvXos8GDQog6w
k5CNfRwKB8PYUyLVEjiN3IWGElG8kWx3/NctzuV1Y2097CnqVdn0tHU8iHP0IdkV/7sFQA0p27Dn
e3aqOG1KxLNGC3rkqCdxagoNIDFkWRjiIazYQYcPSNfVBNXuey9SJV+9BCFIQco5Mjyn1qMp4M/e
vDzKSI4ZK2CQQ/8eRTv6D0VPgPBGnPCCxsdtu+k4trj/itDfGDbYOE2SF27Of3yoFuEQiDYC5ahV
ln7/yfkOM70bQ0pOVB9MJ6bAFWiup2OwodpvJiiGi6QClzpnOi/wpjN3UjmTpsEdonFeSUg5V/sB
8JHDWp1FOWxcIh46QP9cgzXJrXE+T6gnvellP+5MWnLsI64CqXyOspIOlkGZC2+VgVvTVrXcgc53
LCSQDTnDpHru/lrJbYpRRTwh2Wa00UCfXKn0AJbD8V4FwZapkAllxsEBPt5K5HePL7t1woFeQtNr
FmxQhyvhnV1UjIGr0iJSoz0WRIq7Eb+ckA5ZaPufP5oGzRIkC3P9h/OTRrfmVbsxsEuzit9oBxPd
kJU8Jd2ycqOnBXTfyVaNKdBm6JO2sSP9SxC2M5Smh/ffxV8Y53rAFbHq9EiYDBZ63Vvp/+eFj1E+
xecJ9sogBOVptrLMtmg5GNJBXmHAp7b6YMIYlldEgb9tIOfGMJrVP2FXhGyAOrpHGzRWvt8+Uvom
j+M3jl3D1xDGO2t5EH1CHk3fTe5JmkDKcXa4YJVxaG0cHdWlhSa78vUcSIThI47iW/hp9cvwEJci
9MBRNhoYb0ewoxs2pzH+RNHy8ahHn0YNCoPmgU8XejoevFqTVcKhUM+QRD1n8RRh6sfh2aHZZtGB
PZuJOF/Bkvw9U/i1xOOqgb2O22iXMOdAV5zBXYNmTLrOaWQTsbANqq8IsEDmJgmzG3eqC/9Ad9s+
ewpozI8qh3lZNGZxYr17XodLNLRhjVCWqMNmpCufoT1MQhOy2kiddEVZWXOSYOw7ESYwo9LnSy53
iBsepRRrLiYCFQD7/2vSwXD338VHjNi6kv/gRJBmC0bPLRGoEMI56INSawT2V85Qp7Fpy2ZTgfoX
3h4gYevFTyTSAfmSPYVilT0vtA8isVntMzJPbAaGLrxmyFQNlhnPMohaF19RoQeK0yVyAyUy37Mo
fYAZxrOBSne+ff7UqW/WmGRhxNs3fGQh1xqrwpw75MorB0rMMhL2hZHlfVPGpwWN8Egv0onsDD+z
aQy0hTWtRddbe7iGfGhllsy+AHMXUPbgfjSm96ngpIbDkBgT3smd1StwdL2TVuJMowiuPS2wTSEH
7NZZ0p6hc8AADvDM3T+EXVbHVDa+b2kyw0Of38XLPT1IRoY52q3Xfu/tWvP4qvh48VmLGnlI04aJ
P5NBaozA2DDcvh8ydoKiOo2i8QMMSGWRy/ZxdK5jZmuJd4vG3uYeCc4z2EACx02037hTeK+Whxh0
185YLCSopH/ju8hCfILtsf7NguucQjiB09iz6308MuUf3xgJmiVpYFd2aRHA+qJfuEOaJaEPQS3T
LM7eWp/6LbZcjCB5rxY9vFgBrR6kcGKOsFJ5fpA2f+VG3PT9eC7kr62cDtn/O7zPOCnJqZ8Nl/1i
kIyL+gRSvVy/eImsncH4Z0Ax0TaSp1O+8r8pyiKC4MOWvfModPO1q6WGKJDEdqAcOG/kAE1/CDut
tdiFw3tgwCQN/+QGtZrQzujA50YY2RZLrIVArL+fyjST+OreAwin+pgamT0bm7PCaYadGGqvAD/p
l3aZKx8puGVrbHxJ1vWiB9/dQUQQqCOrQPog9K9w5BdEoN9lnY0dhFr9x73JkSEPWl9i+5AB/3d5
Q5Zv2lI8QffKVa1fZ5s+CIOejohnRovF3n3SYjEyOBrAs6yMx5LcJgcM5ULSPGad5uEaH+yzWbre
wklWcwOWeRMTKJZLecoSFUZNLZWrGVC1I4qwcvELIiTGtYy9LLpUvLgpFyYux1cU/h5n0zwsf2rl
1gTer1q29Rve7itrTqOR3gQprZrZAxhPyOS9xVzyOVf6gnDPu3i3cavejwuu8bH506LPiGzVeOTE
mr9Foo10SQWKAS6mHuVPmPBDqvFxbrniu5VLE88ntARfWJiTPEIZrpOrgGo4VRFv1TNFt6KR1NXJ
YeMUeNbStOvfsHsBvwumscbniPcrI3EekoazxtTA2CA1eklbpFapws7CWlrlrvCP0Rjfnpqzo+/o
GIHVVLoCbsANinkQnB8UGxoUJJtP+LK4hVFUhK8/4Hlj1AiN7FFrHDwlBAHbgkX+oZBdN3Fm5X1i
0Mb6fjvp+jeIvhHQuzpL8venBvJ/bPDMMp8kxmZ1PplVzcTmnC8tuZOMv/Me0shtZwhHaXeG0KPk
VK3k61a9nAlmF0s/Ly6x2qslmasOqlP4SPelDjWd94pIDIcG/6e+Z0cNfRvxiHJPifDMSFTUiD5T
2hNypFkpY8EIZLqYHrJIf7Wnb0pH1zzz7as0Nv6Z0az8EFCZcKQSqBouIAKUVas6dC/6saWfsPvu
eIebT/RHYTLXbZL3+sIIQlHQ2ZP4mSDao364EMak2QmiVvUSmhCyWgk6eFAlzbc8yizVqmDeEb0h
PMMSYvaf/F5nO5i41EEtFLOG/sYT+1v2iOi9nySG4s2+W3fvMO/G4WWO52wkXA3RfxguSa4X8Ac2
VzFLZTAW0bwkvbUvGiw67yOw7R6H5a/wTjOC0o4hfwYIDPP1RmMTEAZg2ASGzuIlz++xxyLJREO8
Lm479abADfAR6hAXjA7N3Pd1phlNr1uAk/hVTDkuzK/QA1YaZ927FcO5wOgAM7UXmr3VPbUWTkvC
WJEYWfy2ekxlcdCxW6P6YGxCZd733K23aHFcVI8ZZG4hDKgPb2F7z27Bc8Ypy0kBOzqnK/thKgFF
gThGRO5Y9IvMqO4oXP3K9EUQORT40yNnvvsS/0RLYNsEymElDsPRP/rTYpDoaD+KAW/63dsPXa/X
XGyECf3pz/FXWiSRC8nxQ8ObTOBcE1fbwCVTcDMq2s3eF+fjow7rFVC7yOOqWQEybUYgQS9hRImW
UVdU6K4SoNPtA8S/Tg6OxucZqseRQY/n2G4/t6pye5CEoBkY/B+3L4s825fZ2OvHcOVcmrDz6TD1
5uj17B06yiCJqXA82HpkGanS2OeiS4y0Wy+Ijpgp21wWZec3oNEb/kLHZXijw5asR9OYktc9UPVV
0VKDM4gCdx1Bn6Rdu3PJzlwqo4oY0N/xbTfjJP7EqvyjdjchYSMT/nYMWof8vQVNVH+CSb2SJlOg
WwYR12I3NO3/0dGGBGNMcjma0Y291qASP2uhkuk3yzJD2JyyyGsvSgHwawTayeUgON1zLIElJLea
jnJlICp67dRuMd1u8t2wSMsGW3kqXrqs5t/7GMXXn3VeBK4vUsy/xRLPsBbtVN5N5lJRcIO09bgA
MNHhQT46n8g8bisZdkZFC9E8HMo4cEK/orC2YS7tW1kdo726eprfwKlWSNQTTB5kRXyD4QxSKg7o
nAvJVZxBCS6GaBT5NLGmDwCi+NDeLqIvgkckuWJoHkcg+/1XLuxx/3qYSag1sQSdFhXsIb6OIoBz
T609V06H8WLASZrwxXgIM1IHGcxwDJDi97jt4/WZ+flRYixvocFWNQNunHo4iZ2B+9X+xQFMrUi3
j8vWid2Wn4mQ9ou0AZ/q2hPR6ltaJLbTyEeqTuH+20cDk1x7fpkKvQ5PtrMDOCY9qqsruOwRgiCc
pz9AistVlB24h8vF78v0sy0cPo8PDic/bVjW1J3UoUePG6suHfEGcyGf6ahg+B1d/WBEnPvOW68h
c1QGCmrqu1WyG9DyfwOaiR7jDBoXQiuY5guqY2BHBcBD0uVDQLPkmGavhX7k+o2sfZNxErkcR8bg
/fGY0Y9gaRI2ig+lC9mdUKP76oBYEjR3UgbKHWUr5sJXUZpp02mR9ekc9uLgf+WgeqbsZ/Gm/Wt+
xG+puA7BPnXvVXIOl+1YHTU/SFSc8MNaq8qqcpQ0H3DzCtBt8lWtzA1SShGlrcOgIcaUFqzGQ09W
rBHz63mubCuBh7wy5XvkFcWr0myVcBGQip222EI9+ns+/K36p38+0G4r1uXsFV1lUBo+n5itbPAU
6PxG01FFEOYtC3ONT+nWyFR0K1YPuQhTpHVLk1lFr7JBXnYpm4j77z4n+j2UAncT0C+UPNeKzoyN
dTEJJ3p2byBDOv0u1JRjv5W3HnUq58pxWtd9A38DDnO863k0UhwviBNdMhwcJcP88zy/8MOHAs7Y
2bISuacCMyqdPbVh3HFztghD9g8A2hen6ndsuVtl+Wq29vNhGFsspHff1DTPvdhef1fVyE7c7rKS
7+bOV/GtvDsxGVy7tuLDK/L5mNfXA45y+FYtXl+099ecz7FC97/rPzp0W8yoVrVoDjqWf6TjyPcv
BckyN9iS6yvv08hl+0mp33R3+QiFUPm2W/HSCMNLiGzDKlY6603VL0LxmXLM+Ekf+5YT098mYBbH
8p3n3dIjnLQg9UYqSi0VBAtERuYevB8UCu5s5/Bzyh+fm7iUJibAPgsBM+yKjNHm0see+YKHIKrf
13Is39zn5ZdAHWTxrFZmNdBn3T7Z3dIyGHDbESpcS5VD9kF/Hx4FhlUP+Y5vuTlYJe4Cf0VVCIWC
tLakD7yYwMIwchlc6+cnpHqwW66cdvK5jYu8Z9FyV/jGbFGWDlvp63qGM35+dYOAFpu0F9fNifa+
0BrjQdIC2XPu+OoD0bMWOPFyK/X0kctOrcOBrnruyyOIoCIJAiNDY90KpFwchTBcGPiPLF26R7AC
SaXjKxDFKgWi3SqawB9rI0bqp4C0gMzNHXWWXLMVAB7LZIFL7NYvBV0rimnEd8zQMq3pYn44MVDL
0mU+RoCWoJgzuWKIarBLNGtpO6zRt2OgC7NRqiP35ZSldamTX5wixev3RiP9re+ONCIqplB5G28t
/vjxdGzoG97TszGCNGldiI5EPKUCNwMLtc6doY6wICryL/d0pniGmcuWkx6JiPJSxwBg3toKVv84
PBOjvBGNgotj6UTtiir4tnTj4ZBwd4K6YuNHBtffRu3kEHX1mbk4FfOT31Y/fgkffqkBex1oU9Pi
m5XzM332sF2KyqO+7kRVYEIPFaMS6LRMhKI7sdrXJ8rLhBze01oRIyedVX/ie13srlm1ndQvwwUu
lBLtJ5Pc+xWPDoKEXZFSgUDbudRVSaqy40xepvVQUhKFttvzgGliU2rrWzb2g0a0j+4jq77Vtpmi
8YfOuv+t2qFDgydsQVakJX980MoxxCwAPTokvvBZzVRPxwQJ3M0Y+M9ivicYKWGcJmWkTxAgo5ut
j9rpUo/hk5JdcsDy96//fs1Ab5K5SKYua0H48wYywfw89WmM8xboaaLpZ/Ci5ysCoTXjl29tzpVY
1tBoKtZOhAeYjYkLbTXhiJXt3cBRtD12Goodafkkd2NFlKdxMuHDjK22QmwVp2ZmhRB/08Bvb4L3
9xCKG4Q7Qcuzi1G5ZI7jszlJ4+H/nD2tdM8UIE2XlRH14P3A2bozRHLZYO0RYx8DvvN7xU3XZnKY
V0BjvQOr02X8FNXtoYwULs6tUSq/9QBrMCrZ71ZcszdAo5QyxKbKPiDMW4S9sKjw4KWtsq2ySTaY
kXcybtn/sjs6jpHz/hRXYwdTRY8w3TrUWGEZ3mHRA2TO4b/ccCIvwe9BWHBXAwUbH8q5EZhqUw2u
M2LKj2lJIf3Mdwqnc1fnlQ/Pn1QOgENVQy+8u0ZMcOqGOrl7bjydYO5G5jyskeC2MShZIdv81xgw
ZLRGXYWXkA+RWCOVu58NOS9MS5p1Z3z8AHJwCOhpqxPhSOjzfyQQ7OSM8XRWmM+THz9JZUY4OyhH
vD16eCWg9XwR2ANBADLN9ZDwaEYp8tGITSRhpSiXNeyIj/YmgKZ/g7lt7WXcCnxWHYRXtkRTMVyI
etwWR39FkUJkPoJHSJEeqee1eAYX+JsFvkLwwfm0vWakh9ok8xgyNNf1JPoEWOC/iZl52rw0xokv
1iq79Evh6KzhuDdFB9RRNOGWVLmSWTLe93NwKbZQucMbnVETYbH9WT3uvLDPeXssMQAixn1DPRz0
p9XzP3jfn0odK6NT3nHLiuMaIIeaJAofN0YgjzQKHcmQ/ue8xxNkkS3CfSMAVBXXDUu/c47LzZ86
or70u9V93iFdqje9G3Tn/gLLBt5oBMzmnKNNikVbDk7NlFytbFaRl21scCS0d2civ4DypagPoabV
XuWvcv8riDSViUO96y4FnnckhdpDuLh10k7juI899A8RLgzXwP7lGTk9bCHJHiv8Ucf+hLercQnU
27v7oLNUI9SAE3DcE/BZhHj1Ejg6nVNr/g2kHb0CpAkgs82aIANi6zq3Q7DX2aaONtZkG65vLcPX
YPhr9tAbhNHs/WGD+5Z7lM68X9HBXonvoO3xq9B2vpwZqm3taQaOKf/3zJ0jTm164jb65JVrsx/M
OHmCCSJ6p4EQNLmxKP9qn0o91IrKZdyPUgigvY3u+XcHkPrBorfu7VaSN8ZtEmDOuhfrW/eRcMK7
XEDgUYqlQUcfxTDjyID+OQSrUmVHfR7OMpfevzrFOpN1iocEuMBmXUBYso+DpEXaJZeFOWbRSZ/O
BQuBX5dZbOYGkJpalhHDjfgiEGRfUY+yvO/i1qBtq/6SKraCZXBVnKITPWNCcDX9+JRCDCK1Z3VX
dL33ckTALrSmF9c1CJEZI9+ZklIbcK5jr8eCbNXTKFl3sOBrIupQd/ayzVC2U8A9MXHmOrKUwiW/
fRV32gtUjIu3ENRlIUA5w7pt/XPATcEKONvQ+waKrtPzGTM9cBFeH7NV4tizKFXMCIo2eHfG38PG
N5SymEq5SzblRNMvkheoAZTb20wb3VvZnHvKwolEqZMBz9U2A9F44VxbdRN0U+vXJrL5/Hcv1HvX
vHnw2i8U7fZM8Jso5UYK70tFRvzH/blcWK5yMIWinvo5bXvEgIVIgBb17QzymzJpkUfGLF70bjop
gNdZ5n2cc8XuFmBocZ0VF0MrkBWfS9IogpX/cHvCN+sQfpUz3mmkmVclUvb9Pl2lQ42OGLW20GF3
TD0aMalH6V4oDfzRrgoM5oMYuMgwuv2Rn3sIXXtFNCd2EDGCxMJNubcZfbaV6nd/q5VTNkM8Kb3w
lgq0jHbVnM/cBHO3zpBh7PmtqdU9rMoSOZHZ1pD3nNgRQ5Uar+F4MNj4Wsp61R1yO8xuCWlIfABw
iu/qqwYRTXOVRne/7h500bIcciGo6YkBhZyozf+6sTQNDQAYBMdXbjltfGAR0zTg+NuYeNJ/3Dve
RzYRPgyFUT980D7G5fHucWwr/3Kr94DIxuZLZ+Lj8K9skjpZ682Qx88Jk38cg9QL87NS1b2l6UX+
PR5z6frR36609jLjADOrqPgf43C9bAqJ09RS3XDC09by7E7wKE6TqTsFNy00E27CdhrLfNPWcbbY
2h/QBQsPmasyVl7ISdp+RFNtLGS4SJ3TAvRFNVJwuJ7RlX/Xw6XTskMnqVMhLv1G+c6xEO2NCNdj
qPAQrTHvcgdT0tL8hGqcSnE+iOLVhZWeIdi7teteWr8iy0kpivMYkB4xrwjdTF7nRLm/dUY5O7GP
5QbRRBJNEIB+Cn6ckpHSliUqmi+EEE3DDrzi0c0rxQ6ER3jEciQbjK0R/wthSKSIPtaGCLEMKEEP
2eR5Io9aEfLyuuef4OJo1WySGE6PIwU2qgG/AScQKs8oLugKbUyVoGV4L17Ou2Gon88yfBy23JKI
gkwrhcoj9RfOIwtgEBdg4ydudKstLQdjcHnHgt3kArsuZpRzX3hkQn+nBpV7rwQHgRrN/sHW3jLD
F5YkCIEMhliiRgWrZ9y9+sXBRVYPvfpIebSjF4eXiV7ZGOuG++g6jVigiJzpfSbkAzJA5IABsZPI
2jsJfK7iugsfNjabfAe2DVUe/oOOLLukVcCkq2kGKXzcDnFz2ondjKBhFgOaq+zaK8OrcFsraZBJ
XNGkuDgLwPz4rqvTFJH1Cpa81tIYbYkIece6ylFBoooA/t5iXdrNCatYOhImYe0RcIPNU8TdHdtJ
7U4OiDe0RIrTH9wtcCaZX6iJytIryk8aoS9KIbQFWefxxCVv82l7NALVsO6uNCMf0Zd1eSXPFqQW
VxD9reptCsmN/SRw6sWwK+wVLqQ2MyckETZFpN3tw7tQNoDBF3h6a2g2IQ9nokts22fCCfeQhumY
+v+WHibidTg7nhj6f+C+hXs4osFGvkgLuEbfefjlw3EtscUAkHclWJIKhPGIFFPEZzWfRoadc3vq
dwHp3YEuA3vV6OpqEhnVim2BDyqfk9bonYmYBREOmgadrc1HHl0QN+Y15Md0TnLK1nJrYz6eOcTj
/Tbs/1kAV6FKMA0jpv/tlyf3kog91SGlx/WdI21x2EwY0eoJQjED2cm4UpmO4IE59Ew3qec1bQ0A
DyGhY7fZfSFUpn/ioY/1u074njXdXM1Q/D8M6InkVwgODPyovEcpdlRMWu6wc8XP9iy5VDpKnJI5
2wYBw5Xub/aJIUTuaS7GyAS2aDyfRKYmg1xs0BszEM9/AxnrxO9Wzwl+vQxQh59ROyxoHprUx5ao
0jvUDqZUWKbyBUSFXRfqHL1JWgQc77QfhnQNawLSI5nKtuJxS/KO+guMbVPmF+aBKM3lbHMEsERC
/1z5Zh5SMJZe8BvQ7fNxJWFb7q26A2b40OgeTrRuE1g/2a7hh1SyGx59be4zy36O+Y0YmVSoW2ln
arKyDtTT+NRnLm9fQRFzuSzPf0u0rccGnNa0OMhl52ZJmSjw6Y4k7QQREdKcIj5fMVol2t/CR4Pt
maqsvDQOexAvcdC2c72XS+kK77HrRXE5HL3UZ8bl5wr/BDaKnQK5v7p8J6rRjas0MLyEYCJsufcM
+J4MtxC/X7BjkehRN9e4jnJrv/cJf4jLCTQAbo9JwsdFJEG6gD2kirAy5rLFICbHSMeR+HqUtZYF
Unf2AkXFQH/fqPzWK7xzo5nk9HxtpLXflcwtcGoG5kkdi0nXVNqt3u/xWS4jI8HTdatXw5jVwCEz
YGgSHna9h4q38LRK32bNVPcFQpSM05aEB6MkeVfN+ldLYhQuWMeu7eVIRqL2Wi9czUyiBQKm55KJ
cEAub/NpOkT5oOXJ80FFolApvYINwksYxbiqdvp0HEByZ03AFBvBfboOWUIwFfKtc3MzAO6W96+9
hVJOVDQIfwvKwZlH1lDatQALyL2aTX/5iPoY928mxRo0jbvgTnyJrfOxZGkbRoMkuaRfjnMUpzZr
3WRLvN222WKHGA6sg8o/alEu5wwNBsJh28IThRjkwctEI2p0xMr60Tcv6fMV1M4kMvcd+3QKr2Z9
guctDuQ5S5HQTABvY6uDtH+h3Pd4Zwrrbv/M077lHLqHBJy+QMrLMlAKB8d2vGaLc6OYJC7UqDdG
4DwvmTRyMUHSsOogyZQcH+JqkMQNmrfv4qfssWiaEqKRYlZis0hTpqIBIxipVXSM/YlNOkTFr2Yi
BVXnlp4yyBlXlTvVMWTvWqGfL3xbWwTaTWY1LUR2qfQ9gQXz8ChF7w5POVK+Z3nW+rL0OtfGoH25
WTLkCCvh+Oz4l7z0E03ugZpCUvomOZeiAPcdJEL4Ygoh/jWWZovct0T1OQP6ARErKZBFmQEbu8tX
x1H0170WZjvy8Lu9/0L4D+EK/ClS74xYD667fV8mvMnLVN2WbLbNBnV7d/2cT54OZLvnG8AJis2V
3n/DRd+cUJTcyoM6Km+MepneWHOsKX8VAE7900pV54+mZv/7CLqA7b/G4n3f65/yx3JI+qsfmMKq
f7I3StuEfovzPB3n5SdIi5H+sCNV64y3gGQlWG6P+yJkLg81jk0DoDqaEI1SRYhIESXXEXTNey9E
Ziy5auqyCD2/1UQUUaoousSXKmNk4Ss1PWOi+b0y6EY3XKKSM9Y/XCQK7Yy0nze4f2t7eDQlIKj7
/7KUSzFKxhZu5kLaJlhPtOPsk+S7GkGkuOjxZNe++a48a3gdIk4k8IK33Eu+NiBiUQDsVUF1z4dl
8qX/qqbz1ahiXPIWlwc8n5V+8UVnle34cYLnP+g9/SgS3pnQI+qT/HQu7WMgGNyJZg4Q4/dnLrs1
BvnPKFyoaANEsSacUnIrvDdotfr2l2+3TwAsFZKYwEE2gWRoWmMZPV1afOUSoEr7fYpWtv8LvLoE
WHaOIOwdKSYjLA0LvkBwlagSrZQl1ij1tDAZo26tcnOX3TlQgh2vlEAAb5LQiJ4MQ27SrcbSLswg
NDzVRx6VyIAB/hdEb8AgRY5/mzRxANAgsXvIntIEbqUsYpguV/ydbC6vzcgWfZafsi6HH6rWO13Y
l28kI1P9KQiLsEeKcEuPGQCMwtN7tJ8SwHkjJkkJO+zAT6oLPGbDFGCYw0hgf4bv6ZF1VRfj8SyM
OEWIMptRWU+OZEWqLhsYwtGZ+y19P3DLw+zFPO5J++pGEhdQ8xl7sGhQqPmFkKYVs0SBPSjjVE8H
dOYOZ9PnEIVkgN+h7/RlGDLWxvY4JKVXJ9OEFwde7u0fq6zeaeepLQIeRqOiEwG/5VKkhCFqgsy/
N8a1KcOkW8GeTbjQkplqLiA5QNS2EoKSW87floI/8VOO8gnPke4DoyLIzfXP1HH1qS+7wMa8FofJ
6cGtgQZmuiDoNeJ9/va1qfuwP9dBJ2CJamubim+SU0OluRZJcU2uAJHK9ZXN2Cf9D19mHbsBviyh
rwA4uWK+n6YP0pHp4hyTLLo8/TP562O6LJxU0VCg1eRJ1QoerdO3bAQG87f93kwJBzMqNglnauuJ
WDSx3X9Wvnmrk9i9/OK07HIwlBCv5qPHrZnB1hNL6ACnzDacYLV2f0w/NS9o66IEBKlIsJGRAJM1
mtXsrP+dSY+EbSixzseR7/u4F+50xuNFs9Co20bcNUVfQ086uEkusa1GO7P54EPR9b2yBytqwioQ
pADa9XpcBzQE+DsrNJJNAo1qMNgbMz5ODJec75yU0gkdNMFSySt2N4buEBub/zi2SMQ2jMYNo2+i
5mvc8/v6RxpkBowd0X7KlVuC2qmWVS8m8m7abLbBaPmXOWLl70fxDrtXjg8OuMVMMZ0R2UPtJiDs
RdxiJpYMxL7U8PVr6tDpLHJiK7P5c+4LjZlj2O3M5BP0SdHqpPBW2YJuSxh9q7AjZCsyLI7nyQsW
DsVAuQQoOHRpPXiefyTdPIsTeuR3WFQBS+dKrEc4Iz8YzjzrTCM0hfF5U8+4Vjo7P/pPH7t25blJ
PcFLEYEymfKqnje5QVZkTKxxOjODQMZgs+FCL0EYppKuUzAjFgCpZMo2M+ly9v70jFC79wGDWEjW
qIcwQWeJwg6E7sKdcsPEMrAvZFqQljTvBqqRKK8aALVOxwm/O9BjSFTqVcrEhi6Q6FcrvFHKJ/Wk
24u4HDUlmIfmUO1XuLqRl9eFsS0XPr/akKW9WpLArTxUl1js63D2WXSROdsuyj4v93ATD4Oc/aWl
6DjO8mnqEICGNrS4MgO4Pk1k2hHwvR047cWwS0+RC+iLtqxpAPeh3lUTY19Z48TGjgbQkWqsLNd3
AD3L0tu4A6A4oG6KwJMV7tFUuV02gGrzQJ/9bvVSijJVfVsQb5g8imfBayBpkPPBVfwQGuOhRYel
A+iz38t8gv6ROkPH6Dwvf2K6G1qKxzE09GK1zJnjXnBWRNmSE6Bye4InBckFqYt59+VARJrMn/ek
taUZ7S7HfWjg/OUTRNQ1TSbwdaE3JcnUSSyoXXvn14jSlBNiVobNzSwKVFEZ3Qzn9BaD4NB4i2iG
nH7c/aQhEV5tjg3ivAvBr9HgvsFKsqDJgKqIVTc4RaTf4X++ZVAex1JCVBpcV7b5ZbOy6fonJiyB
FHNBQRZ8s9bQyvwrb0VmEEd8bD+tffsfM+aOEA1DI/IdVtKvSSnKHj2GLCM0bd0hm7T3yg8dw0Qn
hbu372O31NmLww2+cX/sF6flDI9dtPJQCO2eQxOxqAe7+p2uE6q4K8NmeQUTnn7xYLIiP1Ra1rg4
+lThCfw9bBXx78EKMxZ36cPw3KHKp3iJXysr08WKauVHiIHa7bCYcTdXQgfv2DmghmEhEyHSHFkl
ntqAPVf4JeXlQMEBEIzXwUuu83E5I6foDziMtqF4ujylN95RP95ON2xAQjySRDmdE4EhQyhRCnGB
1UL9LVpKXmc4E59JAe2fBxrgUiAClbOc0V9a78XxJxeXJKDAw4OTkDsUNUCIcm6XG8n1UEikVGom
DwAmEW7CEIGHtTxBEaumGKiReCj4mUom585vnl/qk1xHKbwsgc3B/XjnrCdrZAEUzAOmxLWwj3vB
bzKbRQ2QytMXzugXmHE0E+q8C/xlYtXm31Bn7+vl6SLiDPcPyv5sNpjGLx8B/CTSIJ7zuVkzf0gN
axbaukl6ny6EbgHBs6ufMk/eHzgGtTAvtzVi0Ma8Wnxmo7NKmRB/qBprqJXhRpg6LoYeycyX2nek
8+6Sh5oHhP/ni24z/jTuoCqnRAZo6QLYIM/IFl+cngPxYPYxAjvct4CJPbCBnkrvtbUS/nXoAN35
Qm55SEcYowNJNsBEk+WfSZLy0oFzAVX/ryGKsR9c5/B1XQOVNkTWJOc2WT/FJrBRAba31S62BNKy
Kj01AspqoRhjXAE2igYLjtXFzGnKEkEt4bJRhpyCrSKOMKSDpSWrrPz/o2BbwoT9VbJeONU/n1Rm
HBJMtt82dYVYb1UZOabYf4Wl1b98B7z+qhlNXPUIPIxt0l0ZMIE+Pk8BxU8W686jp7q/AuNoIefV
B5Lwnmn0jjRq84ED2T2WmXXeVwzBfvc7BwK7ztQNoWO1i0YZIsAhcC7CdoSr6+EvwYYOaFP6XK/7
Un8+OHzFlS4ncTgnM8AGGgUf9t1RnxP8c8Iag7t1X9rwgx4M3cKuM1itGRzr16IfulBWGVDmgJUi
rgUtgsrhQE2P174Ex/QWxBYUTyDxjcOolFNIA/XXZddRgxQGoVj1oPHM1GuZPvWp16WE1UNZninD
rfpx/eSl+wUHfEiqLz8ZLpDozvDXxOxZwJssO8pMSogHUghL7azB7vwjnEaMMDfMbOYsvowQ+/Wz
CJhqx8kjMkQ7cBEEwmp6lUuRGC7R73xarZ1t9blHRMfEWaa28jbZj2530Fzc5aFqJp3xJDT7VsnQ
hih8lgj4NRuGaJee9byz7gJtJkM2Jgjl94xOhViC4A6hip3wkNk4tLjOiFH4vuuodFHwLxqodQu8
nG7HOwykVGXIDEd6pMFMibblhkQuyRKIvzuXpyXk8ROVJmbMLGHtQqSFl/q6KcINmOxBCzrgcndp
wKdTlvc6ZpBniVAWD6cJ0RJAzCg7imVMo+vhAkCVrvB64RgjoepOBAhtMD/JLAMGZsMTBm/osAdW
9+n/uEPdFlZU48QeoOa9pLJ7ONBEKf2c+eTGK6t7CHtH5wV/G4O1WH9RXX2zwO7/u7v+py5bCLhp
QX8mx2aKdAy/4Oz1dkWYs8OHjZPQqgLTlDHTVPNswqu6jyUxiomr+sXszoOL8uZGeErJdiPjIEZO
r5DXsnZqKsSvvVX4ISVZNrr6JDcNQKUHQrh0k6Y8Z8Oyz47ABaKdF3IS8evIbykMS0TvfxeqxPgM
9m1uK9PBv75vUITaZm/6kHg7msrC9D6EVgmBYF3L6DNhywyisjXGrhjcMCOmUfutxQElqlop0woK
qdq4JNhnJ/37jLxtfjYElR8NegmptB2wr+hHyNiKKiRJ1R3pYH2e2+kNRlHwyGXMbiy3EeD9MhbD
fjF5Liaz0GLITfJrG26awi90CvfTI+v0x0gwXGM4nYZhHKmRRCFU/bPLzcXy2JNWktn3t59bam1V
Mq0p7i6GK+Dq9v61CGB/hKjuAaCq1DRdrursiGyzc3JDw/pqM7Rk2Y/jIU1IuX+iZtpz+KOoJSvb
QaLCpI6M6FP8T02bqzEZD8ea2fANNyhRcz4Hrmt7MYXau1Za9YuHhbLrpgCL2n+INtcaFHazJWn+
t82iEkDrAGYIQcGwYuF9rjUp3QWaHOx848i/O3wn60R7XW+44bCY0YW6hFFklch+uNmS7adnh1MB
I8jeS5rJvKbloXtiAvsm2SwWil7QM1qS9WXjdgNDcu1FZAtjGnqDU2eqAmj/pnKiQ7uw3XW7mCUq
xtnAL/UDB9dvQth/MwRgLlIiuNYaBdpgcN3KGoVUOkFPTfRunbLderMSpMLHpaXiLzQgcyExbVFC
zAbPp8chTbUdE6hiuv2kpzJuYb3QpwcoV5tlRdyfVUIL4S/fic6aWGyFd0IosdmjH8Gau8VQG09W
igEKMh0SjEw5lAK89Z8uyGKOloLYQHX0QJLV3H2gKU6vEtHwHrHglqqkNKBb4Z/9aOBLKmpLD340
Ky8S+zDxhA/2Vos6LZV4iCWV/1thifzJaQX7b8H2hA67uhLa4GpMYNW+st0rbU4otfTxQQQvio9h
eObri7ZvMBB7VJpqRsptzNuNIfCfWG5HSoWbGe/PoIqlLbBRfxKFZ62RuUlXlFVW20nonyvUQSLs
BdTS3BxEYyUeLVpx1+LrjhewmCLDlflvK+YQv9fJ/2skaVe/de+HrN7uLRhaLMBlKLH7W3JrCp8/
/kFu/8A+3uFewdReceHfYBKOKoqMiSWwYl40Nr2c/ZBO4PIIk8wOswZG/tkY2dkIB1gfYaUMuiG3
CNGmx8BFANSmKh6vZeuI8S04ib0hgf3rAHXwtltZQEIn9PtTzsCnO0bwuvQ1tWURW80rH9Pw3Fd+
hQ5Y8rMDtx4v4a1yv62Ngulmf6gsJwX1jx8lZg7dA7yr2MQMhslX7qPYgqtuRPexLLmkMeJYb1QB
+iTTP3ZFeqnRILT6aDUaeKhtUN/GTXSd2MtGuR0YDVS+HjSBgOoH9yeNBnNyPTpS8wGUWtu7XO3Y
uyiA/5hQdqTtjmOzPueTQNUBNvFO3NQM4JZ7dlZoNWVvegs2qwnEg2QvMlsYa3JrEI+nVOs6j2Zv
1RHJ29E5I53Xl7D11c7GTRigXun7kT6d0eFTmK41rQmA+QUv3cRS70IZvzmIs6iMfoOjUzmuznWy
KNlP3O6d2u5cF9aKeo3+4M6F41CpEQHD1xMMAy4mRhiZ7VbOyF4k2rfWJRTvGI0gmSY5Me4vOIXI
d/BCiq5ltrtIv1zZb51dj7UhKjS6PmKzp6ALCsrwgvnia58JZjRZz48opgikA4T0Dfpsx/i4+SBp
v98svyo2bopoEonmc1ycP+U3Bx2MRHKlBj7/A/QfNeVblMHcZ84hN1heOxVKoN/fKfkNteWYoc5B
WBBcTZch2pBx4oC1B+Dh6aPkxOF5Wof7RJ3q2JIRLlJUfRUmXh+IitKdRFqh543eK/td3E2Md0tp
2lmds2IwYD9Rh5M+Ro5ojKzBMv96CWvWn/sxIYqFIEiAqxU2MYRME2/LoAD1+3CRDMPvcU03ZxLm
9Du5S/90CvXSnGgl166X1iILgExg91MShbfxYFyg3rH+5Z379LWLnz/ZcxAMbL/Ns5enSZaFj5v5
z4VIRA7JnznA2nlvJc84U+HnlMQOOqQpzmAhf/Xhm+xNWmojgxSdZ/Bp4RdUUK5d8bT1MdzgTA5/
SxmZMpBgX5meAJBgH+d+D/84QjZ7WH8FdeUJu2BXAiwJ2ub2EDZCQIIwYn5VYb2FHSyNf4B11iP2
TrYyBpoexVOFcO6ueJpzSxdMZUU+UDhLC32aaJvk7XEDYhPWPDTDugBn1Ho0n7bzp/OhmL30SwUz
It35XrseKWcybw2dFAHIuXxibZoXQIrvzTI/2fiAAFW0oTSVnVx40Ypk1lAh39u+Z/zywn72mtML
hlSMdo6IvPKTWwg7i/rl/BK95i+cMAnvhY67yfSHhbpC3Q1J+iWJ3Haj0rOuhO5ytvowwH+HNLcf
TnYUdkCn4yu6c/btFAQxt1cMAQi6GO04pw7mEi+YdoHrO/z55pQLEUaU4AJVKNoGNeB5BZXtq20f
YMyRSJCIUS6FdNSm65k65IfsR20NmMjLgF1vVHfVE9gR5GgfK0zqde/bVKPCQqQSaEryB98O2cEd
EdQYK70aLhGlhUoeoYR/01RrkSbuJanFgWVWdLiaQnO/ZlaVKdSYvLbixT1i+kz+Pn2JEKvesjTL
gH0EglWd6MGLtQuwv5WUPuvyKQQzLIO866DNLyqD4ZeG6te/1FNQdocJ0vdeH/vJw2yAJ3VTpb8u
ZbegNjqF8qasjXTMIIzasTNvrbAycopLHCO5+Dj1zmQ+8q16uuaOX9EPL1LEXvHCeg/8O6VyDx3Z
f8ugWJDVQEgjtOLSzRoDjC8fwR/jME30DaKkTrWSi4MXdrK9qEqCiUNxsLpqntJkjHS37huTRFOu
1mYlwIqmUzVCkhx9x86zD0cv059XuSyF47XGBVsqKvV1LbVJOkTzV8nSiHPYAYXwycFOwRNr+OPD
q/6M+JAJNa7LulJ76hYZTyasLy6trerI4ugaAWunugAV+9GctGv+sANOheQZ285O9+5ZNPidCQw8
sr3Rn9eitdpUKfaO1BrfgFO8lMv7T+gmvMlzwoRrouO7vC9vslK4NAbjeh3Exe33imV42sgnmulA
bIEFODFO6cNsmunfYzIyFcc5jeLjK3C66R35iHJv1bRxoWNmcDHxnHYMIXdb1DyFTtVxDeGVGdlb
s+nii5K+Jh7eK+F8xPE5+AyrNx7eRZ+XcJAEt0N7k+dmLyLaWwNZ2RXghH6iobiYkbSCIujINcm9
T3RQqijl+0dhGR7++SgPR0TuDfqFkfUzHDCJk/Pxy0akYiKTock0fMBSX4nouxMUR14faIcT2JGO
9civdFzJdQq7mQw8lqAhnSBdcBR9T4DZMMlphpQNkptKyWwK3IK3rYm9l5Nxx9CV6PZk86vjd4eU
8Q5+nY4etrL2tq0gw+tlQ7Xcs9i0BemNpbzV4g5AIZlsSh1WX+gOpVaoSbNuAEIElVttQzB4Lf8W
22aekZhrXlxgMSVxhW/15D078ANI3y35de89Iys8YD53uMo1tHPeBqtX5vFu5+RfbZfRx1HTFO29
AltJw1nJ9C+JENp4cpRtFIFfKLi/IyFtw0IU7AUdhkfkClndAkunXg6aGD0MPslEo6KeTJ+Hdz1V
e6x/l/ae4E3EDM7JVZ2lGk/1KoTWFx2hZq1XZhrVoKNJtEu7gP1brk14hQs7Mil3E/ec9/CS/Ilc
uSRoaPtxvjDDxNqBphjSARv0zUyppTGGEuQAo3rPxRpveGLM2NUe9aVrK1mBRk+u9QALYv3Zhkaz
SqiR7hebDreLxEn31JOnpWRpmtMnwlq1Cg4EN+95lsSnj99v+RiWWkej8mJEymmU4siWBDh7Cb7D
3STbva9VWKYep9ZWHXz+B/LHT4+Fl3c5OXmNlCYA+yJ9N4OhHgWg7LoYqueTWPzcTX6uwZvUxXrq
1qFPKdNwoW6752JlSHbD8pqYj6dvzC9Q8MFQKHIcwCE9M5AX4LUPIre/HXEj1uigQgoV1AuIlzc4
QCrSqr/KgDvIa5jQ4J5y5uZQBpyXgLD8BCh+hotrYQ5PYRlfETkWf/mj66MMpWl0pwLJGA3Gz4yW
ZEf5EFS5aWeFcBwP+mxJI7HCYZAPRPjX9Dwm2ZcRtf876ryHvVUey8xLmX9p59k4+Il8RtDz2Vty
WgZMpGS17wSNzvgsd6xSCwWVBqfsDsm7FQi2slIjm7/LUe79PDjXX3K2zLvHU4soYvudphwfJ1DV
B8y5lN/wYpEvJl15dJ8AqW6EtRjUACxVNBZVk+rO5/jfHTPyNcsmIOu/p8s5Ym4vahF2rJLrUZtl
xw+cieC2G77WlaJILBRPkRJHjALBoYfExJV6zTrZgkObg/v+ihBxb5hogDGZO6yaEWzeVMDhMf16
yskQQ6DA2XQAiuG+YyDk33wDSDNnIVIMzPlVG08sXzCq8kg5f9NQ6dLTYYVi8EiHBRvEiZPseynW
lRYe/bm7emC4Bv/RN3exTi6VOjGQ/lcjJ1wHGDBQIz8UYCE2HzuX1ejZ4aN1GvmMOYBdK/zbcD2b
KEeppskrQXGSOZQdCbPvBVUjlEAgY+5BMwC0FFRGOdvzW75rWdSunZaPXNsvxcVgo6xuyjkRElPk
LqXF9nLdndoYUf6TYzVGtihOxFcCwJUKAKnEHeN9DkcMNJt0p1v0uZoBLAa1SpOjya1oxJvINOKu
ns+ti7oxg1zpENGvmAgJG36mg27fC0D3mbFzJFPAUn1kRIEAXwZLk2QLpsGo//mPy0XODKXhnywC
JNJulmj1WqkI7xNYKznenBJV4lK9v9Y/rIA25plZsQViHnGEwVBi2vDEiTe8UInebRwGxhUh3Fkx
TUkOL5jemMV+GPHe37AVmrJrL88vKLU0jH6VIi5vBrgKI5/ty1nJ+QuVorMWWv8XJqhbyNy0I6rg
bCHtMEVvb9WooRETRnRbjPRauY9QjnkARMX0VnY3w1DVU+I0C0Pa49P0Le4fkS2SwX/bVDWVXwD5
yW2+2Eqj2dtzVB6SOmow+8ksvQcjVjqwtJoP7glb5g/mKUOS59poVeo4DZBW5K4OiiSOyhZHGvQB
0MuwuVyeS4Iwu18B1j39Fg5IIivh0i2HXKxkd/UXue+j/I5P1JyVR2lqsN1zGSsBj7mQ4dieP2Ie
64RxI2SFq0H+AEd2vwTXhkB37XMKMo3j7PQ2P/N/jeLu8eVI6Hwa9ZvuYESWxIiE+7fX5DXj///4
Yn6GuzhLcY8DvvwH/tHrbMrljbQlrFKO8Ug8NVuTDuKUg94onfyFd3cFp0t/BhdWTA4p5fKc9DzW
/npG6ihhGx/wHHJdh4LYxcLmx+mkG/QssGGaXQu+1maiSnVTB9BCP3mroLd/H1/FbmOw4KXk5Awz
WYhJlEdCWStxLLgwsYiwEPJzJv1voNET0cHmhacXNNsMIizUrUGQDi4RFWFhJO9Uk3nlYtjXVtV4
iaScC6wKe16brOwqR73uLesAGpveZZxS57/EP0nKlcDnI5qy8CRYmtsIlOmEPVqihzTLCBYgNyuD
xFGP/1rVaF8XG10nAeUEvc/RXySamxF73KJk2KPvgApwVROOEzGOY05tkLkqM6crKS/PNST/G8EN
aMEIGYwlU9Joqe4stIeIRR1YYzW5KAuCadO8gYYUFXleeF04PWXWzGfX2jp6ur5zrjfNIn5/XfUu
iVuwKaPCqIVC1byeZMH0QowYHQoreAm7FbTAXEbLKpENWdXqPenlHC0igOn+oxGaV5ewNAHum1yb
afHG/aO080Zdr+aTYFgOYIu0kCPOpCH3SiS0luLhRVckEkXmQVEN10QCPEqB+zjt8UMO7Brgq9/n
2chsQM9pudfz6mXCZuQ86UJMxwtGek7w8AzcRFN0fjrvXPTHazU3VFGlzQ9FEviG4Si08CS3SF+D
AXm55cwNGk2xNs0TFqtBX5OCJgUgIIZ0yKNtxBGPZ9PdC12B/wQ9wsFP0da07ulCfDkWnKnGY6Nm
5eE2FVUip5Zgguvpw2Eud0Sh/JPgoIVQwOe/Vox4Wu4+eNqrWV5+hbtekXMWsxNH8mAb6WsBcfXj
LYvVTWhZylp65WgwHhEsuOg4mzCN49hXmt23pQA3MfaVye0vcJVka7PwGRiwLHX3IuwqLUfGpPYY
T+ZVz3DWn9/B5PV2coVXnEAoTzcJT3F9nvNZNsvS/kdyxY13ZllNcxxKlq38wMU7vEoVAqzfgKYz
Gxlff0WEzn/5Tg9ukaa4V7ug/NB986uFEkupr4NIBOxnUJuBnvgJyffA9zpusDWfiVxa7cpyZlx5
Qa2jks5ZKmmboAdLWANEwqpQSjdjCgeMF7nZo3o9GzdufmczKgui0/b9Y5BXuCJ0sHvK1aJqk/gx
FW0R+f6syn7P68gYDr+WDkY8BwwBRGVdALupGsEME0qVnt18M9ZQ2/PrrfAS2quLvbKr0PQMERQn
l1Pfr5C55luZ5TdMsszFcnctaXx7ZygPCAE8UTMtqT7dgrz7xhIf43jwGoMdlz6Nx1d1hLBkS1L6
RC6Te57xA/TKyhL6jq/JpO6Y0BbyBg8WvEQRnixYI6DubkhTUiWV6RSNi29fjjaqlf7t4dl/imJ0
bMWYefRUX4GgWLciYLgJkXjmeotjDMqs4QV6CRNUS6B95vxB3Vj/C1qvOVSGytLx1eJkfm/XVyhy
SH1Dg/tQAbI19kWPDoYXzXrLj9qce22pV4pulYdgLrxMNf74ryhteac0PM18LB26Df1DADe3rgw9
er8D8Hkn8GGa21snQ6lNP6qL3O+kwC/g6uW2uieZTdjQKENl4pRUbdlP5kApRxMU9hoqTg7zsY6Y
1/el1b9+0udpj69xiDMsGKww1jgdWYcXp7S50tiD6ikHSe4olwcs6GdwYA2szl/exJ3KijLIUwfY
dT2JrMs7OEdOSLBNFDiJnsQ3cXP3R7d1ZCTCWTVoi1SdrLLa1ylsJ1ABtCMKKoTPYJ/TWIYdP5hw
qVPm7qatYcZ+uszzMMD8x8BnMdZI6Q/Es6UU+UFEBD66lGJMZqV6SshGp5oNwcZ82wgxheniUt97
C4xRlKWB84y99qrkBBoOT/buEY43lRVPH5bHU/NPYKYq9YZ7tzyEJgbVVER1YMg66WdC828oZ8YB
vABikaUaCg0fJVMhaeMLdAezGWjD/Ybe5CpmVWsam4MJ11eohaVqWlwHwU8WigWdc/2hq8a9DcQV
hmDhX6QFtFlUlEcCDEVMK7I/LfSGvx38nPGzxNmkam0MBGr9HHQJw2AR35IliXYFerb8XntsRI7A
K+8N9YLufapEuyf/ur4Gj66LhA3fMqSr47AHqrHvi7mpJalDCHkWe5SPckHH2E3XMnA8cHCK7w77
2VMJkgRaDNW7KIChx7hTzcGoUOUM6Tf0eKb9L9uf7ubMXPPHsQEdJcoAaN22YKkznVCAqa4T9lak
rUWGqqinNYLt0iRscBtmP/WwmzmitbQIsdj6PW8CV0nkp4pMlNMRWXmcaetZwbbn9oaP8iWHgork
q9A1mzjF1uAlaVJjdX+Y8dN9N2r1ZEf2moH6+PTQv4BwktgzPzxXckkm97CLUT5dQI7O86ZOngFS
sKdkQ7lHRh5LeBSLY7rxVuBHx7Gvk6QvzuRr6JS5oye4kh2MwFyN6TwkfgfrQRGAq8A3Sw8KHvi4
EG+89k7J8zAUMWqWJ8JGFv9H32Rd4Wmo/kenKYeq9nfNXWmLzFZngvwxDBUOYyK8RcaJMGIJwU/G
VxI+o3rcHAC9FhaAmInnPNLcxqT8T7GF9i0/atUCpksQgIYp893Lz7gKH7dFEigzkbqLrfvq6m94
GROd/lgSRfvdM7pXwMryEMBj8j2zo7b2/aiwE3BxllKeGL69TmntgDDB6mZi43Zp32mLvncFwyV9
+6csAsWemL5RvF0U0m41DSScoxf7uOz7GjvDBi9cdZwtfQr0I40V7vjR2DMhPb8aCffl6yzu2uRv
puWhtaiZ2AJL05xZMxtRGDOvq0F7tcKG5a5ySQVxPLfVIb9AOvdi2cDeYeAXdGwDIBJBJg3hnxis
a5O0T5MThIoLNJzWaCRp82e6pzlDequSH81IkWrRRlYT5tEIr8wrf1T7agMNEh6AM0oapFn6gXH3
3O2lou93jyh5bUe5dVSHocxe0WkNaYdwGNmpybaHarEFR0RHbfb6Njga//Kd/lMk3YPtHBiAbGIh
sf30EvFY2yWQeht7Xxe+aoz6qlBy+S3RGq/to8hNDBvqC/2XxAehCBkdw4Ghk6KNzBUhHQdrSE2o
nkr1zWo151uQBxAF+rhPV3wxldABur/xIG3PPnksYPkpkdEZWHJa3U/qqDQkT9m43QcqQLW25DCn
0wuqRwNqU9c6uVCcB7CIGWzI8d0TD2KZHXnGiqcRoUZIFsImdHzP9zvvlOpYaXeOzxCM+6wg5DiS
3LR93wPxuzZd5CZiJrrSltQaugpLvpCozKPMUWdWv4gH7MeEP0vSHuCnv2MjjFawjGLaWqm3BX92
2nPmZAymvXqY0ULkMV7vku1LbtJPmtlCmnDj3knEKq/+ZswDZJV6LbxQfzH6Ix73csLTskaAqP8C
smOkRSTxwS3jFufToqO/zRu37PG/AHGwXTNIFKV+tDRTYZBW8lWFT/zNGqWAF9fu9ho0kRC7cd0z
SCWSTY2Qx7ufM64aCmhu0Qcw4hlW3H3og9uN6us+RyLvF/ENZ1ynHzsv+1diuylkWtdzPUosj6ZR
iViyT4oAouIpiv+sgE7cAIwVvpTI9O24yHnriHrrcK7A0mh8zBYc6iQvCrgRdcByXROdkMzGpiek
TgQZjTbSyQsZzM3d8vVW5OgpZQRF8+uF2otVnChSoJQbZhIp3EThx37WRgU7rVrbC2lPnUYplAQJ
nCZT0959grW+FCSgqvlJVMjhAfN/UEAd7XeVxnMAIHzcDvGSgqQ3XITBDbDnMjVKYpDVnosieJu+
Ez3KBMsIGZBTuA6NG0RH8v+Qz5/UcKNAPZeMJAIdc6LixS7PHWkrxFplPZD4Kq6g54Usc1CRhuxA
EDt53IiOS5CwTy5YOQswfviObJ3+gGwSD7yCmgW1A38w3YJ9LsW3bTljUqjUqLKmpArUGmmNqdKU
2ahyRAm0BAXswyyPzzSUt1cA9OT/h4Q9jCxgLP52gHj5YdNSy6Wxxdtiu85LwCMCiWYiSCqXvk9B
USQkn0jEa1stFPcEjh4wEobxw2CTyqDsP4ZVai1kpPVN3xAUGL5prWxnYNGqX9sRFoh2mZVsaJzU
8DuSA9KwI1n48MPkd8iEz2HBVKqEk1nkVQ/UgZb8UztmwDa32CzELjCN+FGsDPL0sq2kOOl6vjiE
b+UFJ/8FQh6mCHV2YdlAAx8qqCsLB0NBV/kZKRdqb1XDz1tUyAvu6v4ffpfN7PY+qullJfKlSeK2
LnikRn1iyH6Fqmw3hnAuO6KJVq+TrwPL8icFCi03Ryt7ZinQrrY4w9MEiCEAWwKjsJBc83b6J6qV
jWxpk1PpJr7uM2nedL4pZkB8WU69Y3bFOYEEabvBg9K7AgzBBUltpmCthQmliEituqG3gx5GNimh
jtrWTv8VKSQ69I3D8BZoq+HVammsnD+5XzKFJ8EL8ks9OFiOcHLaeeLK/8cHX9BvAv3y2owJ6sHS
ryaHB+cO7dgJITd3y/UFuJ30APllESpUr6J45lvNNGsQrt4ZwD6Tye5tvrVABPVuyanAcW7cWErC
g1Z07TOXnabnY3S8+ifv8v8GqKLwTtfqb4blsBmIb+hzwj44uiTnFZ6zgLCiBZGs0MoxMlldDKsF
usQ1wjbb2Vag4eG6G/OzaP4eJ2OjPjlFEoJPoeuTCeyAfTLcCYFaRkLa52pCvy4zNSQRZXesD9tq
P9fKxCpcr2k2CGYdJmW56B6VAFKnbHwwk0sYaZmGdC4nzINZklEt99ky/Akiq8OZ/YKQNqa4Jpsj
MMiAL0vcnbo/XeZCsTvvzoXOM3sjOBFrALMB1qfpMhnsYEFH3uizxZHDauOavUJzqEWLmkW2zzL/
f0zrMkEUIxa7evnwPFMUnLee+/aCVFCa7dnK18BzSnBLCyB1OvnWqHet9d0/U7MPDpx/BlC5uLCi
iuQXELN5qzC7+vw9X0hyMROyM2OkRerlq/bn/4xyneFEOVSWypHsyGqipbZHwgq/h1l9gx9xriaV
/9Cm9ZOe8JMmC47jWyJ9t/DlRT8RW70WdsfOX4J/HXUWFJeBL/lSbxIbDIjLre7awYKzNK1VXTyR
abhhD/5oI31nI9Io9GqIVCbuFVaV5lXxRwvXfGeQ2xtR0QhvhcZCSpDkDq3Q5xQ3vUaaNCBym50P
tTs29wyZVg33tPVJWeOj3ENbmHBW8Rtos0O2pgQK8xATRzY9Hxt5F3mdoouRUb2tXiounstoIjV0
kGb6pvMjw6NRU9EAfViXpCwCkcAbQOkbHx1KHbGbkx4Q7Y+wa4zaIutDmctKI8/ZsddDijHRe7zS
ST8aKfK+lWu1VpL2Ujr5YmFltOT6eA4+ZxuFdR6z6YRTHJilJyNJ9bCiOYifbqk1GJYpSqnmmUsB
IjEs9xUnlUt/Cvf4AVNyaEwbsMygpPkzwzLvNHuuAl5Ck1i81fVuuZUh2gcK9FLSMfX0ceeLpFpn
nz9AlFb9DZbimdjR5ukNoTDTz+0CJJBkH0YGBJez9VDvHe2rRmBYcJqvjk3VfXtxtxNq15OhDF6T
+Ki15u88xqODx8NluLXrxVXEvdo3+4WD2Q+92xZq9PIikK6UuGHoKqs20rOs9rhnlOn0SWGTX1Uk
ddVIgoW1J7JEunpn27+G1z5/6X16TtL/bpJIPcC4+A2bFKdD438XDbBji8IW/QSLLnOaP3jhjurM
KGUPeGdq+zkZ6YBrnKm3YURMYQ61AaHO1Ohbf2xPu34NXww3MiHzewkuf6leigvTuEde/CwsMq0Z
wWsbULGsdWxbM9DTrFmKgjFUfUpyw8IQ2cYi9rXnmrqZUdP1ujqy8jMqmtyRUwX5YKHypaE8imLK
dzFAt65y5LS9scAtfVj8U5deVWeSrZGEwCKWgniJSRlJbLZ8ERuqsUBtvL0TPzM7XM6NjunkWJrm
33OX3PHU/mB31uyS0V6Bl0WgTjMmYxIcs7geG8iIe0+CB3HreBpxhjfncw5hFmh3EsiFSLnxxBhx
mLWYgQcAfLPy71ZMtoIpkmCcx4i8ETLDCdVyupr3KIa+PXTT+4b2nIJUxuMybUI6pHfgRVGTVyn6
B/et/NxcBiB8vkGXyS3o7l8HC/xlfmmXVNd2faWHVBgQNzRCUUO8vN932PTBHEeeRnEjcPDh17vc
syabMWMAky4ffh+Rnr3eCKi11l4DzMbsWtOUgAgQ1ouvtTohBTvzEl3IktW5Rojf0SzvdIoFF2jR
TkfAV00glPgZZzhK9v3hCJsNE3tzC5+vBxGTVKZNVx7Pr4U2GmURNMiLIBLotAIOyg7izXEQfXa4
Z64MtfxK8+VCFUTku1rGboERHCcV7PVR+Uf79w7gwYJLavuzU7wFDAWEArseqfdBQ1BgldCl6oKq
TQ7kLrYcTNz/KiLpVomPEoqnn+tt5mN2UUJmaRU640Dl5lPWGThmPwT6Yo4pvlQZOqOG9ybGhHpb
1rs+9Y2v5cu13IA74ihDW5p1/dFOwR8y5evGBgMNNm+nEb88BFJrrDUDuT8O+ehB5AYkqOBga0Mo
PTo8yG6yb3U7KjRZEEe2iKDF7A3A3Cr/tbGOW/mJ2mZSov0BBQVB/P82i5R3kpNHaAJAbVpAuAUy
mR4fQdI8xY1s49Q6mBq1YMvUc+ziWlruUJSWi3eHFf1uUVM3/EEX3X2iu9p2j3btk5tobaEr6AKt
CEYqQAbxDvJrpR8HHFWQxW5dYvw6r2iELcxArJUXigc8ot5PlBErd8mzUKhQcssw2OEmiQ5Y2iCg
6iekTRI7ME1PmCJbgPqo2ZjtGHvGPye6KssX/swYkBkfkjDncM+/BHGUAa39ocbL6K5ooPYTYHvd
RkIFT5Pkd3mTr2uJ0A+W29m5O/ruqmMnTTmXkwlBVtPCJR7yDvmQ5qrP2uyHCzLna0jnq1EuiJcd
NTtj41ec0dzNflG4Vhmn2bbdZBt9tq0vCwv73ECdfLS1ncHrh7lhpxva1UXiYw1qH91opLq902sG
wEXCYwAUt9Ux88qRcgYF+oWQ8n7sz7vBWQwp35+lRFjWR73x0cYNzSLozgyavnfWDBdzwYrmkN7+
c/EzReO4eJMxdXZQtALKCQ/hudEUiS8SgU0OJBgIMwDuECEF/FhGaOnPHCeQJd4+ajK8c8QooPVX
vLeEVvcO6EMMh+kQvBzcS38GHKBzG6e4BBZ/J0sTgyavULsGw09AkKxGJgM2EMf4ZX+MHANBUA1W
CCvqo/7ZTtVuLQAITG7uGsEguH2ucsw1xTvOYyaxsXyj/7Ke50VIcgN0gTn/E7RHA4Bk1wa8o5aU
whb+zJTXHgcTcBMqwWxnUVVn7sNRzppdjunDfcBE1O3dqvB3ErM2EAiE4WS7kzQJ3pMzeNNUl2eG
xtk6JrbTPJnXHrEU5Ee5BPVmCtYnyRPl8A74JLG+OF6MZ4PUttis9S57FC9PApsvpgM8QsTzf1Cn
ShRLwFavBXxiVYlUNRkADopMpw9qnQ9ioiu74FvmsMMBbkCrHcQHrsPjIktkPHdH1qYv116W/5MY
UjEF9eDBVVF4U7BWf0hzT2ukc3Mmh3P/o9jb4/WKvmDhhTOG+iW5ofkcTlAH0iy0dcP87/2T1Bxd
nJCgyQi9R/1EFHrvZQyC8OoyJeI8fftFQzkQcUtOUe1Iyd0jW6M4lcM6Xw6sYa0Ac9hmNvkSIr21
lMGyhyPxjhbvjTenClPuQN+ZG46KDukz0lq983uJaE2alv47ijnxKq+4525ErdTRyejazROA4UHu
cXp3Z1K2DIY71cutn5SlU/Gx+sPjMkjaWjd8JHdhg5KfreuXN4CAn6aS2otoT6fuWjM92fxK7T9d
dKNUmqYiyAOjIuMW6pQGrhzjU7YrgOL3iq1rpox+Ot9tacNwnHSHxxAoCU2NkzzgP05etpKRIMdP
LPn0kr9mNVlwqVy6DZHKayeRfqriDzZasjtAg2hbXApENwbSSAkNI+ghZ5R/MXm2agV9yOJKiQVg
rYSWkezPPb41aNRX11/JTKgUcj9iEvSVfZ4SJ8s/TJ6HP9lGmzTP4VgnojaJVw3OaR/xLEv8P5wv
jNAti+YjxpHS9sjgCvwwFv2CBkwM2pg8QBN1VKv2rj0/BtSan41I41VHdfG5WuIuJ+zWKIrRGnaM
Gbvsd/fAKR8+aoohrKe9PHBwqmmdwZ1sZXpk8Nai7mPGVHrJhSllmTHI0kYvbvOpeubi7Ck3Rv2H
2QLODEZ15GtdgdKiOTVk1Gvtpnu1xoFhSEsSAxCz0cv9yvMpMnxAKSn5MQlERVYBPD3UhAMjefZ4
38ncCtrycBNK/zvn92TWwfAo6WBL16Ea/KmmavUdik+dpt/CaEEgKWbParQ1JSCUAx5dT7FFqsny
N9mGLS5s1pNkbClqOeEoSApTEIay0giSwQNMpIfjZQLICceTQj4mpxSwWUYLvlyYe0mo099wNOmf
0Ot81CpUMytxsmmHsY+PCrgsZGykUZ9TQ7PAzkD4BprrpLEa9DWmZTaF+Gqxpk4jZ63tYS0OXe5d
s8wKhLbeUjUVP2EMlhCsYl0fEbGvMB8Woxl/mBK1hWQAC72FbnxqVETzMWQ7qiSj0R9FfoCqB+dS
XprYkUJMMN1keENHjm7sLpXoNXkhLO/XpCD0zlHIIbRqKZKVIKTvtej4dayQjQv0LiW6dRmdyQL/
/7+zCT0UwGA2+9+PQlGULFehtTewEG2CBtiauZZYbzePoM07IgPoJw2kEqnkLBxunLIpid0TccfS
lMAuuac1bbooBcyJhN7fWir+3NcVssh1DNpLiuUkPY9JaQAqcOim3n1hsDogEmeKJXLBXd5LeI81
g3aR4TvuWcSHUnZ/CSQlECdqeL7Vb1Ika0W/u/Lmzm6KKTh2LjYtoTIyq+rxqyF4ICKkSe3Xjtb9
mc59OLaJNJclG4nwlybKlWfeqtvlzOF8IOmrnpbJi170RRovviSldc4tL5fjV51zwgALQSsI5OSd
tEe7f4+AdzRH9J4OTv3KS8hZHlhbXeKharttjaxNq3wn7j6aKpqIscpJbeu9RANP3bchpQoCqaDv
fFQ0b+f7Lg9uCBimCnlhXAgnHP5xDpz/xgtN7GQ3n0j7kp1Vj/wfX72ciGaEUSOUTGroduR+FNPQ
Kqe4U9NxzileSEB1Z5SwSOqx2AwX/m6jMqEFmIUSYjWBOGxzcYbfhfI4bylnDJ4Mx58IPYK3nK2A
aGf2Jd4UgsFdJHWY7LhxNVvGiRNNuwemh++96qEmlViIiquoakpJhYGdEHf9F/rqFKjvsvznLqg4
gV6bt3IpkUqNJH7Ln6KwsaTbHHO3ibwDhYGncHYDrBRwfPQ6icuuwJQjlBMjV+tRrWTX5KTr+sc5
j7eBSw1iRDn92v9fpxQUp44sYhsPllpKz/+BwJW/ZNzrMp/4qafjv5xcCRqxmBbkqMrwFRC9B+aI
SRaqRlTf9mXXfwVuFYV9v2RP4QuSjTS+9uk2V1oIfKGzX014P4W1lIUDyfgZP/+TFXjLVk//zt9a
j44o4xdWLzzpaGgP6FBLXuLXY1ZskJqHua/2Jb7G/Ze/TdtaRwgqIjOWD2hrFsVx2qqWkUoaelPm
rktcRnnjN4wstQsnPq3Y2fEjxUZ7kRFCpeFdYICDx776dp17CGHg629sgyvmnLy4peDLOpprTvRs
6XIy7qUNGh2k3YoWd545CL+OqLVP/JdEA2NGv8w+0Oyrr3nElag5Akpt4iy5VLjtDQ1XWP93+fRv
1X7h9dQ7iAWdJaV6yfXZxUi4ygGBAs3TDV4Nz9Sapd7StIWev5r2iovxtm0wX++YFS992i6CeDMt
Xl4hoJ91zPBWeZn7njAGLatr6TaXKob5LxvrldRM59J+lL5iVE9HJ6izxmZz4Qba3wH9G0EA1dmQ
cN7FtbIWyMm9TUKEq0RzmKLPQp+/r7iRZKF5bMDPRYmOPDYgs5QP5oIlLkHrvS4qDFxVMkQCJ494
RuTIP/1VukiHBcwhsHkGhs7mRNj9SLMBP8KT7k1BSobN2iHI/1QdOBzSnWyxXYw2Ss9zBy+erhgU
E3F1RF02TwPJOMTZeNhj8QEPhDtXY9NZqbZ51L3RdeuU2s5IV3OM7itYx6siNnuvodHRcaFOwEV+
EtyggTwbhMHvxEHMQ/Xr+RRZ3CDhYq6QE6NYlvm5xElSySByKKphyuy5XIYCbfdOE2qW2PHIC+zz
Yi6TzX6l5UtVVo0Di0rE1Omb6MlKldldBkuaEd/KILIYTg6NfZtrkmCpTRBfCOZGCVpleqbPkAUb
fgK1hKwDMrpYLUL0bwV6w3Q+4aNixeOslUoUTS083iytv0j5+sBHNXccZekypbvW8LP547x0tdcX
BUTmfYKZfyXrWZAO45XiLcAqXWVppSCw95nEDQx5J4FCJlCnxd9DwvrWp6G6RKLUiIAZDP4kiA3b
Wft8lTewK0AjeeAf6dl3Hr1n9cIpb+pqARw8BV2z6YQM+nlioCJRWdaAynZRduR2lGohJwknrnpD
nteSFoYm68xQF+g+PD7jU3Jv2cV0Ly5feoGh4NdJBTuGsLt3ZlhZ5bXs0lPbzmshtqWcswRY8Z9k
n1Ji0u1ZCXshc0Igk0Hox0WuK327QXbb+J/ti9bwW/cce8Ur92GwErebPDx9uSV6b9c7wwj8/rjh
7+F1bQSycVWTdCQZTjfM1/03SOtq7N05Npl3KuDT5rHrMaGYJ/pN7od6WwdvX5K237OiDvygOfw5
T14E4tzOFiLpSoAFL21QpIO2jBc+9x29m5ieb+HKVtjFJFlDikp6hsVr5bxIf+7qLb7n5KjddbHt
anSTe2frN7e+WerGkAgdeILFG3BVm1JQySlHNlG2Dz8ehEdaCaG7BM35DDY2D0xinNppQZ4h08Ti
bjP6ymwskeqTAh3oJGqas/e5jRdj/lBuZTIYxxJop0SsPhyZM/k7poDyWUynoLRtyAjo+ibtvMnQ
bDP8w5gkMOA+SaxlCwKvmKv1wf7Rz4re1ILS9y/0Il/nOVvFmo3mHbJB/t9p8rCa7JOBxGI1SwRI
a/wNY4GfFi8u47jhTlxOFoYn0WyZO6GxDwBmRljtvhWZUGee4nvMR72JZ4GY6TWrA82YgCBmFQpB
c7KA6Nk3HJJGhH/eIEBYdVbzSal7rkv1HSDcZid85cxtYh5xSE/6L6dCz3W5xEJEHdATfrdpYHKA
W4/Z+gCXODnmMwSYqyN3QVyyWY9kqX2D6CRsZb4XEBQDqN9fifcloSGmG9G+PHSVks0RfXDaG9fc
SJmhsVSOS5hP8zqnTG+hWBc/ncoEVe2I8/iUg6mrGi5S4N7Eyl4B2/MZsD0tIhaY8/IGr1wH3tgK
MYPBk9zUVVTON5prNy1NTA02+I8uBdNnU8T6QDYCsaY7/myUH0eFTvk+o9Thn28zgfzUjq/9LiKp
fkxoO4X8fS2QuW+QQBz+KujfJPzDmZWYhC56154V8FwNRBIjJ+ZS+kY8NTX+7uTYuUuTqnyDqYGe
PudaJVODRMNBUfcC1RZYOtf1OJWBowlSx91WIWhasRXbk/7qMj7WopSXbaY0OlBpS8EOIuZ8EDyn
LXcIKEFfqHxigLM6lJLEmkBiUpteVf1dbaCzoA1lqCiOBRh09JVq2z8rSE0FFaLlSqhYSq6LX3bL
if5vF0sEHpjAd6jIM7i0ngx0rJsaEgPoo4HqJ2S2ldTvXNL6zDyPwvHLL24siw9cYT3C/8ReUDhW
Lm7DJQROdzSavsWrMOPPXRgjikU/Ub+nt4S3Z25MmtOjJYBz9MXzScMTXzLGU9IpiSlDPddoApfo
BzTWfq4V7s0xCQt3NuPK48MfcRbmqCJ51rdsbhIWAUvsGQn8f9A9nxAseB2lmXndor8etbG9i7J5
dP+pRKsfgimiLa3jUdAiEVOMuwjH8kPSyq6RZmZTn2h1DonX3/CL8NtbCxdZM35NtkMjLLGYJ/6c
gV6IJVjmgyVq7Twix0VW4nmvnDCxxMdyCtnpNy3Kdk3YFDDnT5N0W2ZVobfP0Qo6ZfGf2CnzUgfC
i7mR5JE7YzP1ChUN0ycNN9F1uAuRrtXjr/4gESLUgyI+TkG6Em881j/aDNiH/aFScsUGyifHs0MT
47VHGp5Do6FAp7VmSEdgyZpwi/2i7BGAKbrSKX7DbnCnxUQJfHiXPi+TVe9+h/lo9vnlwQjD3KSH
lFdDjxkCJ0w2y274Zep/vircB/kBpVB4KBk3d2amQu3QKO1cgl094/sv6eTmCpfB2OXbFwNXPwl4
pI1jw8Ju35LtdG6pEx66bPxvaB2Jwa8bcx3PriVRBPugo0UV+KGupArGFGNyb2ApPvGNuuRT0GEU
X5uCSoz7LI+9he2FLRyZk16x6xwcN4uWvNBZOsWF+It8JMavCy45yDoKMX8H0Aab4fXQcabizdaH
ogORFtr/dmwfyLOAS3GXhcFOdLYSngmr119ey3rEO+JLK/K0p2119j8BuoxOGA0KTbAE8IEj9oLz
ZbsyQr+ATwdfF9UpPFbeJmaouqsX0qAhrkaZW+y1HtOf1ZS5w6AoYRbjlJbjKCF7pspwnqsGlHzP
wSzT/F1Zz4uYB7ZlYrSkOsKsnJqOaM4p/xeHnPAYUVycIuogdHOuuIp5sAx7bXZ4dIUneuD25ZzL
EkwCxIWynBFiZ3T8ILlfpzSQcUqJDvFGSed3woThUzkvt33LQll7+g0dOVWdJ9kSiL9YUktXCG4A
13IvaJw0Qss+KfAK73kbTE8vAhho9yxyNSjaIqOXcIk8WZC3OcympFnzJm2/O+PraAUQ5yNrrp++
S1yJzBDvEfIodvRvKQtIvPhe3gzVC61gXRSt6v4PRdXrHoicc1Sw78aKt+9znoHne3lby/0D/DMH
Jwbe79Gw5P9OUJLkNqq6XRJHWRPX2TtJJWW60jQN+rQFrSb8djMhuTOa06ipy/ay7nJvrBbqM661
2sqGACk7ubc4Jj62/8BEv82Q4eSrOnWgXuj2/6ouhBsH4dTD2GNH9Sx8FM/0osJABfqiBLE7p8jU
BMHIlfRLKyovSU/q+sEtRd4QAXqJcnRtrks6y0Pdt0crnzr2HTHKZgRm0gInmEEwRuJO7Ca/rJTG
wk4OkAATYFNdpg0MkUPhBw0rvy0DEpHO9He29/xFlsAOp9OjlpzKqfvatbLVs1l+C+h11mXY6hLO
7bO4tmQfvWvCrn4YrxDec8Sam7ksjUfFiDa44/Sh+b5lBHdpc0oL8PTh1E7mXiAOeMlNu/rSfFCQ
0Y9HRX7Ss/oQEdPAM+QoI3eLQyvRVuygfL+QHCMdZMw+L1Y4pi5K2YVsAq8eiMTe8wJZw0COGDxR
VUJY940wnzn5+elYEpAQd0bwEsQ6hASjnwLy5vUa6H0VGldFSKK+2218G9ippCySXil4SKapFLea
IxIDqYsUFysvvDByjsmO4KctXQxzEk590tjydg3MNondRhNQ6SUtUyHJJJ+fLngM+amOlxCb2xnP
f2VSWwS5PVAg7bPo2cN57ZuLbkDhC2ALZcu05UJojjgaqdGcOqp0GMsJWJnP/EToI4KCyuaKNh2Q
QSGPATtDyNeVtiizi0UUicJN1v8X6AsXAtqhjtTHoNoz/zz1tS5yU0AhHN/gXRC5oZtq13DTDw3W
5XB055kuHKXnc/jZ6+tEZlCNOEoZP8XXDs2MRIrErp8e2+k1RvrOh6H3eXp3VhEBhA77Nu+VXh3L
tCwpm+3Y+pnIsNBWRq1GPwJG58g5isoWvaRJhwMBm0MtB6UimATnFifeDmP+HCODih0mtP8M7Rlu
isWjAmnFYSMl+Tj0cM5IxjHbNDjnByIlKgfzH6KLXj7KZ0SKna6Zjrgrr7R7NYyX18GgO1egAbys
c9fD0Z2zC2lNdhb0vRPJED+O8vQhdOwN7uohVT70zygorDndZURWEIg1GteiLO8UTwt2qu8j+/4G
p76FztUjhd9TRCq1r3dVIj50EIAHKkg4cTb3qRRcxQpLSKBxqNazsiAE+puW4/8NifHpIgTGp/Mk
utwWOdiKqIcbqR8KWucEkHPi47132KY0qofHpuAAHuWO/G+G4VVNT1mt64qaRTXGeRxBhQ3xRx8m
SIbPh+SPEl7gJnhCGCCCeOzC9135vavIdWOBlPPEbRx9SUjAzfmNydBxQEJmEWdrTX9nsb9IJaYj
tJ8mh+oDxAV8u+z6xwYpgw7LVvUj/eQZYa22YMJHO32PPlZLtaoREQ2YtWPtYO/VmlQflzBUTUvR
zqh6v4kalCZQP9ZRgr9un3ATn/2Y4La3V9e+hqLqUv61QbAwDXKW0JrN7ne0x7zbdKH1qWIDCI63
OVKuM7SjVprd/dbRgVOw2Hao7FuVHaZclb7ju6AKgSki3Gm1RsIybHc/XHkHv+U5yxIglo9g8luZ
nQdB4Aj10DPcglH4UbBXGj5nvWOYFoZMxYIkrRR9BWZW+DG9VFo+l+ZqrT3cTCZ7EgtDc3B1Trkv
82luiH9DYGQzu/hbulvyXuP6PRScqbbLPUpTBpdxuS2C81yZ8Yb5lNAUubzkpWSVVf6yXiYsGHp8
HLPkYJ21MP5It2ehmLSIoJENyiGf32API42nxh17mn/9mfFwBf4i2HwC85tFj639pTeZWiy11hXC
8l+XJAkE/LOl6Ax1lyoQlwN8tB6VoroHSNzQSknl1nj2yNM+glcfrEIzFO5msfzveqDETghe51rY
DL7EFB7DXzaBUFAzGN38OBZ49ehMEaos2eT7OQqaa4pT4xTV5FJyMBLUPmEbFhFSjhDT7xdT46jW
EjfSul6FfBIJ/mmsj2ASLM+FyAyyqQuc5h6gQgKXTFPLV8xKNouC8UUKZIUJJb+wzS415UlvYXuM
G85MWsW4PL0DHwCummr0y5FLjEoKnOI1GpOiiR/bsacqPBBbVE65noSPS9/udx0O2fOIWtHJfgNq
qq4Mc0A/WNO7R9CM7Tg+D9qKwdjiG99gMKT9Vr5KvOn/1PjS6puUNeWeTsmOEkmQSRdQl8TcvMyl
dB81IJezisZ/MeXHmD7uwfjYpJVebdoWPAdPlaf8hHlZIBv/zBwCJ+fxvOHBf11geDHkPCO+DTCR
eSB8KIWd8TbQ7RzP08O1b7b0OG/C85R6CmAeZAQIDV+KHKIcH31DsZrPt2uW6RsG0+C5GZWIF9OF
RYkoRfI7RpmaxD5gH61N8/r5+/pSjJZUX1Y8XIlTiTBpX9AIQw+x95aPE9iKll1NobLH0HTvYV4+
eO9H6WKrRvOEWjfmLTE1sUZ0T4ecrHumutdZSPWx2OwlLPiKM6c3SA2RSCGcenVMOHODlxNLo3vx
sMMok1Bx+76q0BD8vIhzQL+Wl31c6mivhAwr+PmVeiFo+82/rZvp4qibpq78ckH31t0Lq16Nv/uP
Gli0YMkyT99H5bnTPRWEU8SoZguKEubQQDwcbUd/8Kp4I6LNk8kOkaQ2YmupsC86N8XHLlyl1Cl6
HfReqxp5IWOa2wNKMQ9D4kFAuTIoV0bOH7vmRyTarJ0j0nO1a6mnMToQx0bZ0Viciodq36LZf3vf
t+nfNl1lOzoViOY1TbUKOsxjWdI2DAQoLDQeVGAchMuhUYgcjhMzb3iiTSJLGpq2jDyjCiwIT4HV
mZ6DpTbSPzvSEDacNk751V2UOFUF1lpOljKHlwterral/jUQBRLjclO05MWrDFbXCem71A+rkON0
g3ESOliB7oUa4+l84iedFvP6ONQOk5qouCgRO7/QEeDF2hutK+oZ0XjYh6ux94GymCs46zEXiTkd
y0cAd4lTunsyhu++u5bATki+PctG2i/47301UKVIrFPjKbzkk4gPAFvCZsh7kdPb/54fsiedFNpg
QeDmyRZo+g8/lic0gZtbsUoGGcG54Uc6Ww00fGfCdmu6d3722750AfYxoeKBL5Jis08B+j8s22Uj
/QdEOToL3KNKWjAZpKg+vNA2Y+4UGmlOKSCMooaFRIXBryIWtUVLFkMPEzfgHVUPnAg7jbFTfazn
8VPUooNkrU7OBS7fMBebEwFy5ugqmF5axD51h910f8w9SYWsrnH/wwwzInh6VnkRrKmjbGR2+/9x
QC64Ly5C1OMBDou1XH95vlpOHvX7r9V14Lt/k6lJ3VZb+Lm0g7Q2+RGxd1cEQ7HyW80+3prJXkzZ
ayq24LeJ4x514cN+oEfAAGVKQ7SF2sqa/bfyDS1DOJszWQW0Ct22B9tT/qmbfJ8B7aHK52zUJiMf
5w6Y4M6i+EOvZ09D6UrEWu5zypBw75fBev0rppwLcdp9kC7e9y5ERW6tbkf/jT5hzkfKnDgQJFwK
7aZN/9oLzOZbv+jFVJpo1u9VIVvHp9VYLQ5eDuU1qsYwwAnU+TdwbVwZiPbW/E2iyeanIp7/CoKm
Bk+ihIVNQKNh2wtxxcQd8Vgpjd+6NUANGDta5NySTrobBP8Wdt2FD2Pps7UKjWOIXXPf1gr8eqx/
fSIxd9Zs4xL9Xv9D7Y0i2XC7WzSEt35xCfaRtFKGEIavMoRdPAocDltlnlpG7UDZlxSTXwk1Vwzv
D+BzoeNlKFmlXz7Wa/+nwLflAQKVF9u72X6qoYdXZbKsQRfXzGHckpvSpeO952mYo2SE7FHN9tgH
SS2Lvl2Sqhtl6CHdA1BcYnLq4HrwndLAv4N9kJC86JzSghdMLXhtu0RMkM634izsnV/VP+s1vkRH
DRYHOZWb4XO39G+7yt/c1SYi0fQZdCBR7ZvDIuLXs03rnrPs8TqoQxT+Io3rTspBxL2nWa41QCe7
DH4A45coZXVmIb3j7cLFUhpi66Tmh2cuFqc/eIxBMAzQZMSFCLHVjXvJoW4pYz0BWcbJkPCC5fst
RNzmmSBka90m8rLY21x5HMO6uIdt635HLL7JpIFIx6gOHD8z4X5bVoqhajc5sfr96d83Rql88rYk
wvZWzAJW9iYxg3Jznrt/7NCTR2TuhKaxUuJ+ABhzefKh1Q9gyLGX9wCY5qusoFbtc86QyrLHpqie
IqeN8aRDepAAsxuuOmNnzu5ZLjIBdHVgpGYM2/3YYhXr+YiTgzG1OQI98E244hXGBg0SdOf9mb5Q
Wr7gRoAsFvkVmXw16qFLmRQxSWbYqLAxa2iOrTaz/H9RVNn2MMms2dxS+DptbsropyAdJBFTA36H
r//cbf5FK0abO1UNuJTejHyauNijP3KmcS0EXjIP6T8rbxI3Z4Ntl0VjA9AL2RPYhbIgmXrV6cI2
BFux34eABmTbdh/yU0gP5j3j8xoh1bBkfITMjzs0q6b8ZSGyxZUoHZ+TVOePKzXO0CZ82yRO4Pny
Z0MJWP5pvtnC7ZaFhnjy4bYdF1FRE/v8S8I8Q5cqbQm0GxwVuMYwXASnovbHINJ5339EtOFcbt1P
MaVMHv7QJlpu5JEW91littK2Hozlf6SurmwMQLKVWbCV/wK52ijOAQGnSnfV38eWv0x2cTBI7XQe
+lYx7CN4MZseYFreeeoa9PVvttBVS8cymXLP+er9OpliGMCYrBSDKwHjghGOvUcMYTX4XIQA8vMi
+/WruDWCwm9Nrk5AezzidJnlpz6mk8VsDPkuehnbd72uB1df0N6bjYPcqanVMifL3TIyPlFSXaJ7
SO0C83R75XoIb6sBm5keIOcTJtxEeZ+xAWqOrIvB2OJWTqqRgKfDAKoHagMVkXZPgxl140XsES7i
nnuemVQkATCaef4CdQV0R5wXp73rCR9lMPi3+bsdglZZopz8FieU4A2adRnFRtgxky9JjlUzAVe+
T5XkLIRXLdeWyOoPjWMfn2rouXK2p7/Oct/NI2MQLww2RgKRwdX+eNqfBIIoh0gXQVCYmiCl820w
NYKsMVz8Hstj2h+9pvFcMx6SuspDGXhW/8qNh9VaucA+HPRSGcAdPFpeukh14FSkF/hE2L0MWMff
MqNAmsZPPzmYL9JPrf+yADr3qAEFQgosoNoRrYsh1IpV4IBF+eFBGKPbi5l0Gj770BoFmrG0NMlo
TX+e9ZUJOK0Ny84z/ZY/N7CK/bWonu+n8L1uGSwEHAHDujSOIvVHWUUF/fKJxd6fnCi2r9CBFzHd
IgcFt3CqR3U5BKfTG5qGXra8isKUypSYGVaaPGwFSaFEkkjMdErgZpy2V5I9uVNAuRsyCIvwvC8p
5WVGIRE0n4DlzdOQcdhJbJn1AGO6SSPo4lfUsv+MoorIX4utFjRgrtqgJ/7HX8CQjyaXkWmXq616
Jy4MOO+0NUkXeIGOJIRgn3W/cjGGIXSUs51uwv3jxr5sZaKkByT0aonJD5drzJwHWCALANXfF1tz
++PSMRQUFSKgmgFzYoqFN5TIoE35boUpuN8ykRUGPYXr4aBXr3aK9tvzAJ15Nm4uA7heWRSekXJm
a6iKwLS6J+qXm2sVjt5tTnlc0p7XBmKffZC/ELK8usU5WdT12Z/AyUYK760RxeWdQmj5n+rX3Tze
GGC+kfkKpBoLOpwgrUigNC5f692ufv1vxYJV3de00uLTbtPlYSfll8ajb1kr4OkDg1YrcAvxWw7n
BX9cYlljFnHKE8JcYya7cKd4viCXD0ua1gRuYJT4Oe1GnHHDp/OaFXdDHgZe8yr0raosn64khZ+V
h7wFWgEgB76hgfCElqgTQJNAcoUMviEhgnP+Wg6I1CTbyvYOGe7uEodpJDK7ZdpUVocPXPmpb/Zb
4JSDCUN+SWHF2Y/8r5gLGv0+jPHhHn/XF8+uS58Fmfc5IoN8CFDRI+wNKRALzRGtCpsiQcq/HDcY
Lqm9fOxmJ0n0kc89VGQNy6HzP5CBZ0Hb5+DdjXA8R2XQTBfA1hTHODXI31UEb6lSZfURbM1wo4jG
rBxb7cPNlbRJBLAASQMtBi6NI/bABEmbWeO/EXV0bMMV5ZLW/LLjXJjok9GCoon3tGiIhup8DA0z
AlOGPrhZryPT9Xod89dTByLa7HLgmOrUlkgnfKPkyWBhOV4safdEHklDdxHK95nNFT73dl3Hr/zr
CQGNyc4DNQsNu6A+T2nMFztcHrSQet8k/E8XLvuVmtGy5P+ru6upYBcHEXGCjsaEdCckAZqzKtb8
FBuG4oA+hbEIy2Pz5Gcqn2mLuQmEivKS4g9rdYG/bphnwSeOrPKpU0u7T8A30bpowHcrokAon0ud
/I9n0n0CMsid0lLoAefZaO74+q0rFveVIm34SUH9rjCg1wSzWduBaw3KaOhmx/OcdKi089Os9dM0
I5E12qZS/9s9T2rNri9s0OM9Z5nCcthiUpuUCcTagfzwi+OROnjrR/cY9GbPmHhXNkUv4kYThYqD
EwYc5PSEsQnXc/nqYOhdKua7hSqcnl6cWaeI9iwsvjya5jzUBR7qto/w7bc1iuYRKmTWUgtdh4Mr
9eD5YtQdIsjy3YGh16FVp748LE+VJuze4jIb9QX7uQYO5PrTUPVtSRW0PbmFzWjI0nzQiZFgV6+k
O7XfPJ4HrglKyysZfJXPU8TdR0j4vbaetF3/Xdx8Oo6WpHwJnqYiq84eaTyt3Y8PJqIbn98BmZi8
PfVDDCbzo2tA2v2gq2fFTy43PDGqTsNZqWxMk9lhBIL92b8p40oIlfd6p55N165aF953QZqWd1O5
GZppaHG+yin+23784C7YXKlKJ0kZg5VgAHyVkO8lTT4wA1Qc/nrHRAfaTyG4nhABx5NlYaD0Q7na
+utm6O4ChvFFmWlAurMqSUllgSz+FGrG1zU38N2il1PhW1yD9XtYm3RA+MOz8xExLILnoDtPbiAQ
tSUfz/3WDssnSHFtDhVIS4d+BlgKkxP9OSmWIS/6QIZly43FFssIKsCJFBm4bjXukmxUyFye3/X1
BtCPxMUIMH+DZ6+/oG9vvI8bRHuRrGbhgRgGwgPL7+xjEdEck/Dfnfg6IhZoAySaqQj1MYZS/Gdo
yuAWwFgFhwamaSZzzk6mpUdd5S0X1IEhhdLXbEN0q5JS8mPv93FrlItM9Lb0q0dUS7K+Y7/7ULXU
4DjoC3aDtVKmTr4nVWRspsf8dVuanZ8iVRh8G/pvgTe70TCTwVX4Eecr0/TrMREU/esThI75DW2i
9MJwuUE4SKRDe2rPWlY5Dp0P884X8tqnZkfYswDgBCy9xcw16QNCFdysvYf0a4tRmckEycv6mwX3
FV74NPt9d0wLi/ZLLZlvBx01nqBDzAr+97ZvqzxLzx1ZhoRRhqbXgUd1d7qijO+QSNcJIEWLyxob
XsiqQGvfJCHU3BHWDvghFPZaPyjA3PRdAhsjV4W7+gM0hFyKEX6glIRZ5TuFDgA2y/KaNhah316x
cJxZkXdQAnjdGcjqP8ZZEZku0W9cE2xa/2rknu01ybFLweXxk7FprCZ02QNKTHZG6nTXVjY8qzqP
eKFGB3lyz7MyrAohBgd78maRINOTLZbY+xaelwfYyarlaU/MiZUyL5BLbSJlzZfiEzsOMIsGB3/S
giIBWg1wbspS7Iof7+Uat6BItnZkLKbuPBjmuqZx7L9RgJE6k1n8SCOZrAopjBNqGI85soNoWNCs
u75EsJZCqcKrzR4/J0yZfA/J7tiKK61uUKvCYoS1gWCaqU065/kpsz0eilNR4pr2TE2FcjjQOp0q
K/U14EMqGo6Ga70bZGU/syoh7YqRRyXdOKN2If0hnpeWPACC0qt/Pa5wTaxwpQqgwVAE0jtCVbFu
mEgD17s0niMiAzKKMa0es9UXcGY9aMR5YZhHv3PA8KUg/+MKtngGqjFgHR7phOF6TuC3C/h3yZzF
bEB5VWSXj0QEPKmCGVTb/whgv9Sp2SEVxcCaaAFbSYB+/s7f7IVIMtTvwkuyGnghtS4MZ4+72r/c
77sejpNbNLfHHeAuyqXl5GUJmsKCUAXCxqWVGcy9s9qxdxfWYZOp0lcvJm+jywN+TAw2xdxolM3Y
NyOOXNY1eaRjxjSQaIXaBnfbOyvnVg6LZN0Pzd6PnhV4t1S+kMGG5QSDYXKW+wrJCINy0HRqvHur
RtyW+UhambUhJmfOK2mrXqmRE8bPDWB4pkO4jXe4OttzyVCcYmVQk3f13+l/Ov4V0IwyvowFm2Mg
V7p5IqFmECTmgp5IM+VLoG43ctOvJU6/k56JLOONkJyMPE7GDjYr6K8ZONyfBuJ8e7A59U3XEJXL
iMTLxL40hF2jL1gDIW1BZwUbT836NqYvKmhR5bfTDcyFXzea2oMkxpZuVVYbgGsPSpApJUXQNLRj
CMCAyJngPLp+58xqd+m7GFuWMOwx+0DCvMdam0niK71k8bVmyUeyCmlPiGfIWzEN7nwsb4xlXLhh
zELE2a/Rh59u1Z3CQLp7jUn/o7Jyfi8qiGio/5EF9lsXPpcXQyCklCOo3hOBs1QsaDnXb5VJIrfo
Bd8LLq5ifh606DfK1FwFOiVq9XuCNNLaKkbxEoEVMM+mGeW1z6d+/w/JyHjXhzbr+xsXipa52Seb
S//rd81FkBSt8d8IOt9qOXkn3QiZvGaBWj83tRvbdOAKVizHGaQsdm0SpOS85o2RSrToZlOI8qEc
0xpqqKIhV1h67W1Ry4UHdKe+eFYwCvBfbVTUVuOhYetLMWBovuNpWsj3+xZztHAWPk22DttM0C4E
2LiAS/QnDEOVgt4iKmz169uzMGTg9VtRCXwKK/JPxkivG1Naa/tX+gAaQwLkevlNf3a5InurIzUF
jsE6+M1dpNkKSSmPY1fNDle9/LmZ0UMpHwyGHFx96wKmcHD13ckPAipxH2Msj0SDzl4x75WYzcsM
6PZQarjcNn9cw3PWdxU5Rk8yLL3wnYlVYZZ4ZJkow9q/dilqN45ty4RIeCvJIeOVHTGuhUh9YiKw
0nRV2cK2Lu+Fj8zRszB1Ef3nWSz3fbOsog1iFVj5KXSuuiA4+D+RKm2AMVj5fnpM695uEMq0/Yaq
OeFytBBo0GXJiFbykAKwv53sHPC2EKI4tFrQyqO1MEk29MlpGcn18hJlJgi6kB7/MCEdeCz48Ci4
QLSNt+DXdXwS/p0yZgsYy1LYm1mIwOS/MKWFyj5W5OQS+krf7RClR6XGQJ95eXCV2Nb+rZqfwWQd
/nFzuoEWyjvJJAhryPKj3e0rO1WxGztLsaLa98x5a7XGV+B87QRXWJdJFqaObJE0poebNA1QO9GI
BAc5y5HgRJ9Vj1Qemr+rUwfWZYPHTiQfIMzhKMqgvS+8YEhpGyCAs5eUkDpW+ByqrY2DKKzYO7qB
BQPBVN9GgpZrcsAQZHntkq3Ei/h2l2a5Y+gaLTAUe4dig1i3Xgi5T++dssxFEKdOIiYjS8OShCE1
j2JlLYkZJRHC6lwuZnqg7UIZSr1+1+iPPVpHp0lXkKTEJx/Mt11NOxGB5y2FommCMQiqPaWsOdnO
XVwFOYjXpTq2ZjCNjoYgzkT6PwhwCQSlQukWyW2ezevx7o1usnGp5aogty1kzvLKZl+sMzuInqhm
EzixguF7G/5gSj7d5w6yelJW3LNG2WnLWfCSOjh/Vs9QDWYk/O9XDriTdByyxAFIyF7IpWXHVaQN
OgYxvmjEni7ZZAktqS/i+gAadsHozKALNdYZk+cYDsAIMzn8YxiiC1bIFLqPYba8I7/f5WQLan1A
wpsaaHVVFEAsS9dmUGVlr38hGEeFbkd7ZENlwslVGq6HHP4ZCW9L7ZowI9XWyDYrDfpiq/kgNPLE
ISfloQauzgE/EXdBmG4K0Vd9GtBLnFpv2H8h2U37a1AvpWScCs6fhkgtqQtXPzZpfVnK2byQNoV0
tPHprQgpGMIw7Cy1rnVY7lup3v2Lv1rvZwEXTw1xOjFrtMuRd0RydTsyw6a4bSSyzAp+K36bRNjj
F4MBcgQfl68E2/uK8cczuLbZN6UQp/3GvZlXi7Ln1LN92sJtLxeGKAlRSbahSrnAJK2XqCnU2UVC
d8Y1qdlSdwsls1fx4LlXmVm+LL4zTK+eANqhU5zd5EMFxiTbfJZI3hwvAgi9Xu8YBv8YSvxeyiP9
lA7ZW2LsFjB/xezbFP71sGEHhAtMtyfCheeFT/Y7o7fQwYWGgRwfEXzOvRu+LkbSlkiIZF3t9efJ
911a/1eiU0yiu9FJmVMFPDGHLGH2QbmZlgAEO9ROw1F3lMk5LVFxGd8Rjn968tbDDhe/prxPVhE7
gyAywJpymR0fdKmpQVqiwKMWS68BpySVbWAbeHIKsdZES2cAusuoYm+Fs+C+hGoeVDgrXwQzTKCx
hbV41YL0Ad49OfH3dk0k6Fjalkz2MOLD9oFaLyYq+ZfUItsGfF1jShmhQ2nBBlXdVwKi6n25RGPl
tEh9XvWykx4lWVFeiDP4aZ2TCgzBxk97yOf85rkLTDnCdXow9MN9dUJD7U3UeXOqkhAQ3lF9e0gf
nvC+sWgh/r/DtJ8loWrIRzs3xE/bIRGkErtNdAJ7FufolOCQ48UCE2gscU4uTH+MWTtXnqPHGbtI
km7wDkQVkWtWrDtk2AXn3OeJiBVVRBRyV8ik/BAi1tUP3hjXHDGqGW1lU6qw9QenopsSEAYWi6mf
Sj1LK9GRFGniF59PPDb5W6NheYLW/O7gtzpyoq+/b8sRr0rLgJ5h83AhedFirnK2CAptj7706sY6
zPh6N3hWhx9VYYaTOY6uGEX7a9bJTh4T1W4SqkgfJ1m/LeRJHMrk2aCLW+P8deSEP8Y3lpdOYzHE
nOjgnlrfWYQ+WR7z3mTp9JGEt2Lu2Jfzy78g1xM9cfVDkmMN7jHk/t2kH7cxucs8vk7tqXHLyHME
5PeY4HOMVWmJmFqBbe9AbuDi4cP/ppaS97izTMAWDDLodFcp5sccb8cc/6KYTn+4uLfxEV1D9R3z
hhYSt5e2eK2p7X04bcG3ZZMVF0zU0YUGwZXC3tg8MCCLIFoT8o9Xaz8xuE5kGj0nSh9HTt2QCYIF
pKufuQke2GDA38ULhIZN+sfHffjrFMN1BD+umk/n01dCdBwARQNgu5T7DAmnJjI++QOGOH4ZP1P2
c5HFHwqY7a0bQ2Z6DVq3bMX2uioNU+rbs//9YHsyXmm+SXjw+5UFcodsFFx3je8W8jD9U70pifIQ
yvPhWT5XjH0pU/lp4SOxRJb5uIzGIQlRND7SF+Zb0nlKjjNJW257CsxaCPgddNyUHcameJFJn9qb
9HAllmfg0Ybv0krG78CnMr5XuZjEqbOrm7XSJfalsbvvVclw+JfE72AyGbVyTpocdXu9oP0FfyZm
odFz10HvSX9UN/O+Da2P8lmow3lDeW/YCOzpAYn1Z2R185KTE6nVmFa+vSPoPtaKudyznXU86Ntb
9C+iauGgSpDGK5pbGKScAcu6Xd4lHovzT74yEZtISCmz9IR5TqnvJ+kl+uNt1dQpdsdTJd1Esz8F
prhFG5CVMNYUVH+iV2BQ3RUGTDfVUY8z1ghzF7nLnaffaPicbCRUPYzvC7XtUI+v90lFZ5dNqfEi
fmNPdtCi4yim+AWsVqnS6SrFuXt37QGB79jdGINLW9rNJ9vhohc9DvW5t4QNoz42Suv/+Ezk7VOh
jrk1iqJo19pnMJex0icFh82WBI491ITDmviDYv1OVLl629elCYBqAUXBfE9fNORcbuHiq79xu3h3
MlxhGGS2QR5i3o/1Fuc6OqfCdt5gxpRbOoq+3iXqyLBpZjo4bfY4YlFGEwKnvChlgWNFNyrnI9NA
YN4S3ucAiHOWXfDT7qh3NMahUy1Eckata+KNSZvTTflNHhPAmraSV6q6mo95EzrHD7vt/uMYFR3I
bUCCsFuSISbaxQK7pLVl9pGQMFJ3wos6Vw+Ii3cNR+7s00kwI66Ryna2A/K4hxF+amGnmlbYGs9q
gyAbBCVJ3iV59ZUimn7naxiPrVB2M3PkNU+oEtkkmGOFc46BYfwuK05V4C4DA/sOlk/wIj8trThF
19yMJ19BZ3K1w60DhKdxCC4Z/pKBlfQCcpYUYFfyC7PJe/MjzVy0VYxt1v92RyZCo++EZP3iq4iZ
QdLhJk6DMovUGI5/nvdakWh51fYb0i/8Rp/SkW1nakJRitNwMqdtydD5RggXyPvfijJnTyGUVIzr
voDKdkFBmyCEIb2B6qVyrywniUqF/lIlCYarU+q9gMyRR/X7z1EFtjp1dQiE+RIoZ/XBnYiyMfDI
xjPqLpK/IBiAH85q4wEDVwzdyzCAzx5RDQdUMKYV9AP3qsrQ6PC4QLB5Rfkex7Y55ZztxI7wnITn
RU6sDUTn/y1uqvKCxhdGO0u+WpPootXaERkdSL/+oIMfAouPQZRH7kes7EX2twCNGU3oMVsSmdSe
oaoP7WYQuJx1XFrfF+VVgRdHn8kfNGPnKfWj1eIlAbDlmR0z1oOGSNtBAecaM16d1sZdPZ5cCo5N
o3RA7P4XO30XQ6yVfjpsaWnZ17+nXMLHJVzrZVXWyKdCxYwstIziWrlwIdE9lpG8yPS+i3s+eIQ5
60PbdW61oKsUXsfrpJwh8CclLw80Pz2/370YxsCOL73qocxBNsMXCF2t8EiGsNf2rsCNv9J5XP88
DHSAKkEr4YJsLMOZBs4EQpYpJZdHyC2jpkyVouk/fJjDd28aW9VNvxQlEWgnYZesQphHtORRh0be
1NlazG0ghBNbbUo0x8twbLmgLUusOjFJ0qIsPKKlIjYewYkDrxvKNBPV8tBnEs+43Yc6DhYGziV2
9X7ss6k4r0IopWS8wTrVIkEMRFo4rWd3L4B5LdC06fGZY6pIsh4KF3oZYY22bSMMhaa3rfKpbkFW
B4+0ofHDf7PePDAQaeWryF0VrviafksjCSXmorcub7ikGwucxuJqGbXAkZP9k5JQ2ck22yhj1+PG
vMS7f6ztDN+Hiqh6oujs5sNhaf4I+QrY5alYqj8ZS0NLnxYKDhjAzjMdUU0uDCQRHYgsWM30d/XR
TDb+SXuOftfo9vPzsauSC/NpiKUMv6nR2UeXfSo7GMDfy0NEUvkEUW4/6Lz9VkPcfs/hpUBNrZSf
ptxbtYerJjKx3iv/SnIFaVvS3JUeOLLgiL6ZOjspgKP+XnN6pN7uSsA4z3spTzgdwtqOykMQjA2x
N9V48fQ6x71tWHCKr1v8UfRu75Kv6CfchlUEOawDXjg8gzZl9fs+wpLTinMBwQeMH6kgtti+via6
2smaiTRpbi82DNIKcX/oR03LFL0paRMBulIORcpDPhhxVcqkGwYn6EhRRQvOgDarSjHOG+uc7CSn
C5EOlX/jTd1JPfSTetuAgLsXpbnl85KWtxsWlRZv6Sh00GlBEIXSB8KaWl6il85cBnv38dT9duEO
Xnv60dwHYei38UWr4QBq+/keDWOWWjn0TIA52z9N5spnuhs5661S8fOoR8GzDrFl4qKbeRKHyp78
bjd5Xhz6fPGPbPAZVikHeCiZIGolYhXXWhcMP4VkFPISeZaOxnFXCunbRuT7rx2ucQG5t+Pg0o43
AGCTwFtRYH9SsIsXJU5Jc7+h+j56nLp7b9n7xyv6icvTyW15P9wqJeLxH8TeP09PFV9y97irJ5FV
WLQjHtLYKVBb5fwpzzyioIkT+94cKfO7UqzKSjPwzd0m/vW5gA/9ISzIQZkqhRco8yfmXwBqavRv
PsEAPPF2asCb67azvM8lkwcav//zdwFIeav/vol/wki6KI+nl5C/SCk4M+Yq6N7xZoiKyrlPcJA6
nSqHwIK8Xo8bAbeE4cSqSaIuNxwloGbnx920SvTUnnyOS6wsUiKAcsddj0KByUFqWoJDfbpbtrkW
K0IyWozWMnqE9f9T70WCTYRL0V6j6+IhuAS+AXI3O945D3VR/T1H48hWo0K+YdRaVVGP0CJFNuKi
UNf4/dBEUo4Ts0UyS50y+/G7taMswt+x2cjy7xeK0WLkE1L4SU2d0XLWhtAh+Q48TmWzTkLs41qs
4GBjBg1bwd0NILZzXPG21ESHg4ErR9C/jsVOgTmseaTStC0WdjwmHWvEylUrNeTN4mDgGjf6fb3m
YTXjqi9R2rmFCEI0ZZVWCH2jPPoFmJ1SNV4O1t3H8wmXPARqihGwYA1sqF07Gn2vJSUDIqswGXqC
fSxLuD3uKxPtpNG+U/A4OwoCPndx7z1gt0zFDLSkFJjRW0Z3ZX0sdqUfACOQWxaybYHtimVk0uI6
IuVmrKyGoapYjt1ZH57SkrZC6OENL7IL4heREBAu0SCVajllYe5jtunQJkiLdBHdUNwglbjTJokA
TnjxFvqvhfj+1rqphFZZ09kKtpqBcJ+kCJZr++86dCTBVlPEz9aubu73Y2w7FG4eavpGYA1i/Ycr
nj7uD4HG8s6DECvCgVTmbx32l3AHnU8UyqO8dJD/lKoUQ5wfBkjpu9AOhTJJFlenV1wrg9oVuJnu
GnmZPAzZ1F3hVMnbvVkf3ydFay/M9oR0/JGNVOn27yv/P6rSOoT6JWdgwH3oNMHNhYygg4cxQ3u0
dTHfXv+qksJ+VO+O6rQwpX+aT0llRbfy5Fp3KqWIe7ldXmemHqQ6HRvl75bpa/jfrXtk35twUkbX
3WBkO9GdS/twzoWgLlQZD3IjSyvc2yCTll2XSuPrSXzrqTBjq9UBaD+9aAOQ91aoC+DQRYECExX0
xDyy2+8qRmlT1NS5WSkCBgu0LybWHxm8njJgPrpkmQG7FYaUlddFf58gxI9lvuVon4qo41tazs0L
WjLNG309YHowN87Er7LYvVDMeeaGphxFjOsBckD5q/UOOBk2749ZE2mtYl7r20glyRt448uvzMjH
LhKa34gYF95mtNfNHVLmin2IeC730pEFALC/oisl7GvO+LqVF649q3doJySTHBRW8cZUgsM1porc
olBTF20JpFABA7jvJYYOpcaiwUgCTnuHupa23+NE5sZjxK1VlJyJVhuvrA8RdSE00JO+2g+oTlDu
71jPG/HKTBvyFwWHEOrbw5qWO+FMlLnHlv+/52o9I5WP9lqZVv9PmCrYrc9ANAWjifrBx2uHoG7T
CreNX/txQA032O0rCkQYI1lFEg14g549+Dr//S14NhtNn/i1GIyWKD16vfS0YhN1oqpSFyQ7OXQ7
J7jU696zChx5lEceHbKPc+EsKztg7qJAREE1VY8iNQQF1BK4bs66HB1xkt3oi8Xpud1NF7tzI36v
oYOclnwia+AK/EKKJor34Zly06YxaJO+ijpMPnkP2lhvB3q4akEvZn112RaEmwd5skxsXaZCgEyi
m9J15C8BAxIMY40SBXZUZRFX8IVorIyIypofIAggqcwQoYt7zufmC481WnOccu6VzCM9VvBCHh9I
zQbhOWjwjDlkfr9VHx3RA5eWIpcnBVde6tAwPYVofEaiRdGilqoecysBNwX4lIGMYW7WyaNZsq6N
BkTdgjnDbBvWMGay3Oe6S9Fy87RfpG6UIu3KqwB8uhZv+WTmebBL9MxDA0j/Wj0gkHZvRQJg0BeG
fJi2G/pH1vqoUj/+0lyOigDP2+IHUPUhfctNmvc2WRWxjOrFlqk/faHXLExS9bgiVbh9LKrxB3iL
jKfd9bAz4D3MHOBNRmP1I/LVK96N29714dX8aEeDECBgPoVUYUgoa82CJMFfaS+9yLgZfKR1Okzq
BbUaoS8TD2itWaBQVGkGSlv1+aO1q/uWg2Cq0TCxR18uRvX5o6UVQnKr4QDGZLPUlUZKVZ4B7gYO
kTAl6iWQgrNOdiZapezRyj252sLe+LR/P3yEwe9Wa9drH+C/KUOwJGCdBVF2zi1G5JAW5mZNzFoD
+ZAF6BtNvU+V2EZvVn25bi2U+HZBI9M5G/Ln/UoxiN9dfOqNn9fWFkKSLZ1vJZ6lNx5Z4l2Unq8X
tqKLm6QAGdo3GtbouMUwOwNw/Z+mqGs5pRTi7aVq67dvgbEm+KBSRe15n7WE09zZTAAcfAO2wP2t
2cCgLNfr1Q/nUIoHx0Q/1W5EuP6qBCI/zeCXILG0yP6gN8X2kmFBfoWyeTuTXk/abjbrQs4MqcHp
qOdizCZx1BPfBBNFfSPjdS1LON2PyIROPxcM5pt52xOmNZ0Y3qagiXzQoqZto3JlcAVRRWuXXUQM
GmCqmfrEc1cfUtqdn88dP8Y7LDhU7Ctie1gUU84EHsTkM02oj33vcvbfAJ3Rz2bB1/eha+/6frRP
gzbZ3trXFbhkTSS/6+k7qNIfNJ+6JYIVatG5DjIq7OBAeJEfaBYCZkYl8qTlaKBPHRcB31gH8lq8
Du3sR/3USjYvGqYFI2jPd1Wzhb+JG6N9nHaUS9aIz8I4+0Q0ANag+1GhZhH+Ctl3o58TMXpJXgS+
HXhlqaGmBthsVB+Rdt9jsHTBEkxcVkvp5dfWp7DRr/WhRQfMbWUpvwdHcKVILTj3OCEGU3rQ2M6z
Rvc2s5JSSnKid9B0AGhQr+H2KeIrLJWiBHeSJkfR5KuTPOM0J9YXkYtyVqhLoS9qoEv1JAIBQmPd
L42doDgEa5pHC3fZSDm7/CJiEi4UxU7dpNRkQWxS5FUouzc+E8YLZi4TIqXJP3iCKRMBavI818vk
1KDaplRx+iz6CgYSFHqLMRmC9JeCz53OcuGvpCKHM+v/qxPyPh1SrUqyJxoXwWwfQ5QRR6XCL4Z4
Ty45TUHW1JHvKrJxcSBdfewzm+BqQLnbp+/m0PvO8c0O9qUzSy2V0N7HU3eS+1XbVok3Av/iZL7N
s968KQrjwmdC8e3gZyiyCLfxTmD22Rsm7QygnJt/jsUIsB3kG6iaVAEEVGXTAEh879xBMWQwWuoC
Ui1OXk5yj71lFKZerXmM6Xh0/tt8QS+P6NsazxFCWvhtjxF+A2Ipvs8b/mZRr6SazXrW3IUrQhSo
bzEqwLPsnYTLDVAEdzEKctczr7OZqF7X7MCIGqbZmHBHlI8fnPRIcrmoeJLKd6DUlqlnTfRdfLdo
5pWgartZFmGkcWmLJdCQ6iD1SMFiUAdx1EQJw0NkHbTDHLOp6c4Tjcggo4iW7/v6Xz3FVpdBl3WE
WbWud/34J0b6sl2cUeYZPwpNbX1bfRZWQYkys+0vtg4FaK4Zn/THdC53ec140nTG2cFVPnBsJamA
arjEUQg0ktRQMEVP631JGttUdPUrQ5FfFsV0JAJPCU7/nDiv5oEQNc1QYl/pHhTMgTyLJV/i1hoV
WpgjakfHsnw1+HQ8LXAcR+fmJydZb+pi9+B/uRAJ0nDpZAUq3J9syorGG2qJKbuVwTkpctTczlpH
fMKWoRKzQyXHHhUbLQ8TwKIUVTmq/szU6OxPS5gzSyRHxTWeJAYkn5ewceGEadBPzsGgpOttBNBL
yOzZtawgNnfymOA37ILZ+W6B8PbraxisT2vNARAF2j3C78ITaK9/hmamLTPSLxZorjMZzD83IISv
iVdSgMZ7HrXqWAoV4urSKBLQ6upBwuFRVHj0RYiVJbQUIUM4U2A9Lnntya10R4nWzFaddPhDYja+
PD/wpktWxhvwq7uRFVfg/L3FNgjayx3tv84pvza6YGjD+lXq+XuRl9Wvsm0VWoTNUHjgVrDs2B8o
wire9bEnthMyeV8ptgHxgY+KHVEDB3ygLwuenRdi0d372twqb58P8sSMZVWKlX6vgE5geKkAX51R
MC+XFM+BLn5LyExB2B+pMaGsKK9/4H6TaqERFRXrHDUjmvIcK0mmBofUEl7+9kbkkFw2otRuzUil
Ht2g752QAGJyKK/Jk2ttw4pUOJ9IQPoD8I9SALOgMug8zgKolxFhJY52xg8zTxM/qJMMMazUXOMM
pQcPtuqf/3Smk87fDw7Crfsoax0MvgwxAfMEIswP2fK2eevvqZGNKyBTBonK5Sk9+X6w1S08yQO/
OcfBP1r7VvIV93JCLGHfmPhU/xOwI0MiqEZZZO94CAlBPG4+ALS2smErj7C6fYVA1vBxHdsLSw5E
CeNzqrduBsc86k7qkQlss1Flb4Fq/naJYp0LvmfkFVu5/8EHt1IHwl933USrkXFG2z0JEUNhKg7w
5qSsr7Z4bqleo/GiMiSk3i3orCSsmdE9LlKHNoUiICsqB1yGfWLHrnW+0PlqQBB/hmxNb+zq8Jwz
1qZWP5XCNqBSHYJzmn1znDvN694SgKlgyQ1BX4ftBOdbprcGSWdFOK1aFihNfg68T+0+IkkA+GGx
LUs15JC1G2c/WPjZDhiMC5Nl87kmZjJinMZLaXap8XusKN0Duaqx84oMSq1REQORAT15tevU1svI
YI20jGCDuvq7aKoPAAlj9m70kiczOKvIVtXJ0ju9155dIVoVJdCzDvOtiHGTXFduXLQgo550T9nG
Mh5Jd1ndfr5iha6F70IpVlrg8AtmYLqenku2EjTMuzEVYGlCioxBc8IrrzI1sCCqn2+AnP+ElbUr
txgmdz9dOK3IuRgRdls510QYaFaxnlQ9qVstV9uZvUrrKljA53L4g20Vv7+ka7iRxa48c1qHajRQ
3oq50hxEgxwM8AEEVn+Z4UAnqLPwaAAsz4WXJ9OGjexNJZpH97TvhNAI+/LthGbIc/jluFjSd/IX
Gi6tj+B37samROMvwgDly5vP+Vbb8uOT1NRaqXb/nHH7VEEz62y7YZQpsBFGXmiJ56JcDizb3Mhb
3Xk4NgviYGp9ktd+sqnROP/Cmgikwalton2jQsao5N4AokdtwpBd80I3gRRIjxZg7yVkLaAj5LXD
FCNlMur8fG57QqkSXJjJe5wxACN5+YxynBwbH5fyVAyCscAyejkYzPOo+IUdGLJmJhSXrM6+72i9
th6liUrfKqTfSXymNZKsEoy2EThltYUeZj9RrscRepflyoU+fnoYa+fJnjvhGUp2Mjcc6GVlIq/Q
1wSXdifaR6e9xnbrRgLHzr6b7Hs3MyTCO31tgOZrVdRJ5Hg5AZoMK6A1FSVyfG4EdyaOoxaVYmgw
RuAO70eLx7SwILpXYKe6rNTLKL0el1t1lM3tAjAgO1jrEW/5pqa4PGugMe8gX8UNpCUxKhEMthvK
CsitrseX/N3DIi8VX/2ua4XMK258BrCJ50vht3Qb979SUpCXqjbB+0hWdGaVqOl85F/1G2p8ISfP
9tle3A9Temor6r6VhBWFAzmQopi9Fet1OVUYQPjSVX80OudJOSvamXSCrphcp+17lXEwqGFxPCLx
tJNCql3EoJgIyq9GkVPUgGD+zjmZhSg5nAP5tx1F/xf/x3v+mDNSjjQgN1Xa3O8S+LCdbF9p/qmi
8cqQ3bzXWfRX7V/A8pnXu5A/HNM4vhwj1xdwf869Y4aEG7+m8gye0Y9UYjswfFAw42AXoc2TASnB
jSxTev1P7UwpX4tQBBXD0w0XDL9Me66/5J0wlE0oN1JInUpZ2b+VudG6rDKC12IhM0jX07jVA8mA
+bBbkxbKmSDKq5MEeaSt09JvnrIlH93oPlhNCIktbdRxMP+rpD28ahQ60KAV/WI1b4CCw89rAw4u
k0gPlWKDdQDyPLG16TtfQJs5f3GpjGqCuIvQ05X2BIPoiEvYdVb7E4vwQKRFX6LeIY/2AHYl7NJE
qzaF4ImxZwVP/9vjkzxMywhQ59Rr8kgvfQJM+4wk77LU8jpgj0UWcQS1CFH0/xN3NCQOSHE/yOPN
M6UYyL6SGiTdV5OnoXiEglRT7/r+LkgIO0iEIW18vdSYVlWvMI6Kp6ymALGC3+2kFbA5SQ71DzGB
0vHasO8J0cxUWKhqUQmMPrXIrSrVaO9K81M0xjsoltqU26w1M4H7B4eKn3cKZqWy+lZMjE+IaEH+
7R/TUHzVeCx9WxkIM4AQQhUkmZ0+UQgJjp0JImI9Zn59dgY7WOmODQSc0ZhcCQYkUtkCs1RJwyom
eMdHehDySxC3EQnrcjWsXHUqvqJ7W51A87pI4cL6osl0MALqBxIYH/SFO1pkv+apF2lutA+AoTVy
kYVvkQoONEj5xVVPPX1/6Cw2uJY75vfiYrZO++b0CP+uuRdJVozvXWrxIut1JOeGc7WSNQYcsi6L
1GhExGTuc1ZDgVq/fdg+4XSlUE2lDA/4E3Ea7tptRzMAujmCmjYMv3tb7t/nQW5on+tOO46sjG38
wsAAsPPwe1B+04o1DgjQxZm/NVprkm2Oa/p40+fKnBQZGYec0iBf/8dmpIz2ppEC0/GyaB+4UKW+
Cn097Rdw6fkVq/MjnHidm/jfvN66dWXqye37zTtTNzP1mzaV2KQZ3lizQWF81WWzXfQAxmVL+idn
/qay2I8FaaPQZxCPJ6SAdr76FZPEmbOv6HZUf4dQvqRHYyZhR9OUBUcDfHho9x65JcP6aPOoWA+/
MYZO2P8+NDb8cXBORbMPjOFiS5FY6mD0Z89aD1XXpObzV4w6Vo77emWgdLvf3kXRP97l9tPMBfFI
EWtayFQuWshHGULy8dnVCM7zvpf4V0VZzvlxtn1ZkKxLVzw0WzmGFzWhWFy20L5en2r9+z7iFUvr
CCUP7Kn9Q8NRyHvsAWcaay82+CvsAElxrpSsCIK06WLP+/ll3qC9Fal7owE7CvFc6qkc2vJmhvkE
CdQ6heIHObw8lJvV+oz6KGKbCZwWx5nH9O5hKIgXYS9B6uz/sa5tWTuG+eg1fTiqyl4dS2tcbPQL
Qy1X3V7K5Gsxzkg9VNFPF6ftwh2u/0JEJZWe99j5u6Onf7CRsrDQdEwYr7zSd2VEEraxOvbilxxj
bkV4dEWskuPd9DClLKLyNuEMkW5ZGiKsqHZS7v2o53afhPlM0V3OkCcj5/5+Jz3GRTdSJ4ajpJek
FLy5APxY+hnuzkyuDIvX6UGhHQmuUCvdWDe9ua7W+25odEHTLv+RHcIRwWyOXcjE7gb11E5jUlEV
siYqr7TsDc1JgdL58ZSslEg4iD1DfMmMliMbQl6jPvn8o48NqkPoPX8PKuU6UT/elQunki6ZTIXu
6ogIuBxsynUmTodxB6b5xKEDBLlL6CYU/5RPrlbZjqS9NSb0A26QPUfrcDBZ52SJThvp6actwz+5
X/yWOYgLMK3zEQC9jZeT8vt/jRSmrIqngE0W4jA4uj3CLKTPJTEyiXShyGvDzThTfz3lCmXz/sMf
WKk9TnnMyE5W1uePU5dL6fZ8IlURvswbANKX79+SoFCq6srhq+cCUDwsP1SbYUlF5SP4YD1YQMOY
BYlocIY3KYqYttbPRekRvx4IeeOO2TNpPS0hj45M855mmphTlJM/ne+FSZiNS6DYk0yl83+13ot9
CbW2rlvvTHepJv6DvAqFP46ksf/GeJNEWCnuiikxHrM3CEfyjpiCZweitjWM71dI4jpmlfePLF/j
pmUxTOUlvsS8mtMlBnaC27SKj4I0dSmqXgfAx/lNSVXYnIDEwUOGXRKcp+u+Che/Lk9hg9qRGjYj
xfGWWqU7hcc/tjaLCpyh9FNXIZcR6fnzHgpF+c0UHivcmINYdBGP29BYICJ4pfgeY6S/jjpTWLuk
JXfXDuwIUkz29X6veh0uk96wi8X2iq6LU1MrNxV/jlZTfAzsRx/eIH+WkU3ieFm7HTelruuO4bUo
ArjOQV+6wMefa2hbmW1r+ywr84ZnmMZYLCU6c/wIfGZF/R7Lv88sYZO5/U8VySWnAwwYzVDjift9
Bz10grlBCUgjaPIMiDs1MCjIyfs7BWw+SbilomjBPQyqUMkox/AQOZQqFweRpodVYoVSGgzmyUfE
bDU/VeFdaUIV8LHcJs63/6kNYPjUwSyhvwHfZeEeqH1CihC81WR+v4ReUFITnq+BDd9i9NK6t51c
KuYb90J1bP0hndhxGmJNhVPJpp2+Hu19PwEB7blxJyLQ5oEilGINPKlRIAicIlRxWcRZIDDNkN4z
wmNpGNxK/2la9SEsUgxqkjaKAUjaKvu6y3gpxbNXyq7Ofa70+NzFhTZs9NEqXg+8RPFMD4FoEcvX
6pKeZyL/jwHzx0bbd3ABjYiuxMi5nqhCW45FwvMjMqHpff27yxct28erTawDVkzyVJ4t22ye3f0n
aYLUxDUIZFFVTyBRGkEiwFa003KpKVW4KwTOOabhF1kSufNqceUzA3SYlckPVxJpdKJq3sk5cl9N
m2zU/Yad+0ZG6Ay+7f7UHSenIcmeDSwRWkLMDVg3yywNYTlrqNzrZY64Jwe77FIixNQLzTNDh6UP
Rl+pEIDa828WZzuCanZES7FUQ43gCzMlvBPGhInz5n46VkUaIA+ASsqlDQtYioe9ubge2I6/rjyi
FRRagtf8aL3b4gCevmQtEuL6iHFzecm7rD/mw+DlZ1FMCWEvDJCoOgdhkOMUDe+M1PpZNfuPmZlg
Z/ChPukI4g6jjAmaIg7iJa2GhnjCnagMQGUFPgNgdAjw0Fe0bF1HONosXReTwOUr+18QN7cssz6b
FWl95mugu5WKAm3rH2Sp7nGqkz9iEoOwM7+vWQg6i8XHVBbpoG4Il7r95EJVryJRzovTnr4kcZwO
15lJhP3oOKLgMjakxYKjVNxGVYzvDpnb2OCEEt16nQQa2d0j8C2tIQN66h0bNnG/T0PFSvNR1Sjg
dqDYmuPxumzxQjtbnz+cc4SVHW1mjqpHPqk9lJb2MFCwCP8ZgiAlwyqR4XB6lQl3QrK0ZCH51m6i
SXRRVYCIiAwzGC7XmxOno4cLwKz3y64rowg297M8rsuoHtVasVr+iEcu6APnkmcKoWNOHpf79qCI
u0iR0/0/xbCbcjq8pBNtsc1/vAV6UMDLGgq0bdJpd8xPbkB5iGlQdE88nQaCYD6K+hv9H7Pbc0ww
URLhPlAr8buqiMJGz3+p79b9UiQgS9G1+cQiAPekZAjXvcWhKXC7M8erNZQFEsAjvUHBpVzB68lh
36wEpazkvbz06ebBvNKgPOQA/rQb04ie93SBnlarDJEtCvaknJxRVGT6AGdphmXUsln9G3aagZBK
hChwmEjWIbz5EVLfn0zI0w88HqwRguh+B7/mWq/gTSOjtPLREGK2tX8C+RqbqnY8yHTNfww37yw1
s+FMtIcKVXZfgFibDFOUcQX+Af+Q+CkYckH8/MgpDKXbFETmU/wAJWY/F+zUjMWIM5H5dTEv4/7o
c9il6+/7WHMTH8VQHZvDGcJQQVOvRkaOt+dmvcWzAlDlkbBdmzIZ2M8foQRfBEpMFKzZyHT/WJJa
YmiEbQRKablcul9Zf6Icgsr9VllMtHzN5BP37PkRg/BR79A91vXLc0ZCyBwjfNr30KMiYRy3rXTN
PzH8XpkNZUS3zwEgYUr9yxQu8AYRqXlCUmsCkS0OZ0xKW0o/JtNHnGAXcoufbUj3Go3QUVdvxVYh
KyoOa7NcMCFJRxHduYIhRcx0EstZx/wWHMI8yy+nH2HqtqDGJWAX4Er4fLn6zmQz3HaYuvudeHFX
bVjCL6gbg26/89g06MEG2fd6FGnJrYMi0+aHn/vBT5C0fyVGOBxslkbD6F9rgx+9qc6dxzn3TrAT
qYCmz3F+8rXEBWvjljnGihaVs203PvAmIAQmrlsN7Z34kZnUJetTa5tlFop5tRhiPxoD0nlOWvyI
2SX98EWMneJ+HDHU4tT16daFDzA6Cfwcq13XWVDdquwbcUz4duz3EdSE57XaJX/+oMLKe7PwvgWz
qSMZgsP3d3oHZDBrg46P7sBE0lMrbphImm3jpZvCl/OlIRz451xg4BZTsGf3eTt3jgklbAzo6Iou
huMdakMK9sztSyIxhVTAKBNGh6NunsUZod98akmtXRh2k7sal9dcxOnkwXu69lYidgxXEZyZ9OPF
JqFKQClBy/2qWQ/lqVjzbpW3A3APEfljkib8xbRs+lVQSRELipLpTu+e9+u1zGvaViE6xYPPw04O
OaGtZEl7CirGPGAkM4rteedmVfWBpoMKQL0Xxx/GyCcWYIBbZMiiRZRpExTs19GcL8Y8fNCHnY8S
ZEV2vvb+lYsE2DmasJAIK5de4K/c/nDcdnrxwl+7WkmnNyaNazGfXYBs6N8WygSjkeJBda1kp+U5
F391FdNueQYdqDGzKoqSZe1GgYp6dUlxiHnPYXwfuvDIAjbD0EkSElSP+cWzOTymJE0RwNcoymVN
BXHqoTb0TTtdJxgcrHmEpzsUfVjx+uA2TIa20dXNkRODJ5pFQqNzTNQLSgiO9ryXbHncnh7vgFER
gxdTsMz/NPBT/euc7DuCY/yiLqcatr3ADzuZF3g8pkL+lX/DgX7yDjuX3Ex9+z/ge9v+vb8XdNlx
Mdr5wraLbDWU3hcxJJYBZW2n+jCmiTB0eispel+zazrQ3QqWz5fX+XUycKNsroz5Gr5VnlyFZ1EF
nRqOIWliqF0zSoRxik44ysjdglWxF3YeSX+PLSXdrBYvTR2QqsKBxr4S77DFXZ1GGyTGkQCY6qHr
UQgwmooyO+gohMHKQEgHfvCOo1aRvZQDTbH8/8QyyMu79bGe84Qd5goxSc2wX7zXUDtJy40bIFhW
hoxdbZimKTUArC9C3snLzCd68YVDeGi4kZQmyeQgCTMXgWLkPVfLMd+qY7aFpHZIss8icFeS/+4F
DFNYQGJGqSqLzQQZ4tXQWTobBVr1ex97BHMU/etQW+TJ7EyIdjjxqOOLPFfFqX9CE0Agv1dP2Jes
c1p1pdskDSpZLxr4w563rB2yJy6QwLSeeSJH0bLReW5aV4Ddpk+dn+mvwniuOdMMTCEoId12IZ6F
uVtXqbExDX+rzROVqk1cbW4+db41dgMeDgrpC8j5Afyht3JN/L24nSNUNDpK2upxbffNiAdLiX4a
T0IPdw/moJa9tcxG8eypgYTOEQkWea8ugKszue+zMK/xa0EJ/dmV50xkjpDE2PMQvek87wGzMVg9
j3BpydQe6Gvds55YA20SF7MJOyg3R6dBBpWF/0fkXz7+ZJ0BqbZrh3t3Nn9lNuVpFLaU1LyU6axJ
7iJRQjfVv08HiYIYzwgPCZKlrZexVh2srqiYApAY0Q3UiI/XXbfUpNdgFX5Lv9tb4DeqDXXfX2vX
Ue/QiwYRXKysPjmn+llfKd3c1zcpLu065Ywp9wAKz+d0jB8cqnYP3WhHG/djizHnl/++KNeZMSDb
V8byUnh3aDTtoeNnkAHowh4n3z6j8Z8GtX0KiN/WNBnnobT59j3/HYHBCDPgr2cobj3Pv95olgWs
U95w7ZAgUmpPbKMKmxDZGiXFsLJ4BUjN7/+9AYh+K9LYsI/rSaFuOWx060z4BLs1SeP4asRaHQ0j
1pu87c+dBmvNRcRjjZVQ18HazSPs2iCuMZCM5LRkpnyXPfUkMRLXoPtOV2UmgNUn8ZAwZaXjbbky
BO1qFg5/OtF7kb8XVfi2NGlRQX2niCT1ADua6F5mLAQvi1io1UwEWqtLEfyZMYTtpcMpC7msrikr
ILO50OxTOTAH/A2V3L6wwI6yG2R7Vfyw/BJVaiadYIY4oZxLacsl5PBbduLp3c/zJBloBdBiXyHb
EKYp0Qu1LgqcxPBuEZpDyISF5wnF/LgJMSYmu9BY0eOXSddqr6c4SFIG0vufnDgs7QtL7rS8lxP7
rTR5hwJ2S10Q0FVUt/wtimuYyjKuGTWLEcj/UOe2/p4clTMSOwh9623FCJcGtGEhv9Fwt+MiIGr/
y2MDWPVLHLALB9DwaJpAW3ZijsMgkwZp4jY2L0bvXeTQJAEqHt+JHpBWR7dOIO5GrMcTC21lTM6F
jK6xoOBoPn3GefAWHxzwDr9AVpEjAAdZvNhZ1ymQNqIJL9HnxNSSODFTpWSZj5zqfgDkyJc0u/8r
CCo0Udj/bBR9VNYZsPWSF/fXhNMwxTeSAFnp+z0WJ+PZRvGlFaS4vZMiFMT6RdUfHA25J7VPYSV4
ZR3voFwMT3SORezfPK0V9uT2yRWKeDGCsjZQLs19fIoIcIrHJ1UNyzIUiP0soi6FsYHPWYZox89g
u2h7zItIR/H+5bJgW9Vh3M0B7W1pBakhm62Zwht+pf+RbamYgeeCq2rDH8IwZ2VI9m0yN+u9MdDa
ncg/DNlvDHx+0JZmXCCP/HOVpMrioeA66J/B+86zjkHcrOJKjNc5MwUh86hnE48TjTzjBZueFpW2
tGk5W8N+yGQcxKJ4mDNHPnNLl1P6YVZ0YuLmrql2G6clMPfQ0D/75EdMevFcnbhAScMzHueX4cB/
BXctsUzxRO/rfWP5ZdUGGfTQYzQOgNqmvUlaUCQc/qRl0Lsa64zTqGt0qLCsKpOmUv2x/rLMQBBt
FceRIDOjh440MMP97LSCnl55SwEC/Xx+9CSV+11GWY/iJJx8TJFdmETqUCv71T38leaQT8x/dp12
X7m9jSeoLyCJsMzmH0ztRZflzxsx5L4ePgh6snqjYA5u4yEHzioo9FDpqBG6HgSa9iLWxpyTPQIh
54TqRxMCs9FfaJiYvU0j312rRjtd6flIPL8M1qwFdfeHHF0gEMlvqodBTBioB2TiUmCPN3lxTKNf
dTqIh5qkb/cq1x2NtBQDBdi18ZJ/W6fymGw7FVBIw3ZpCu/bw5Eyg698kl9RJHwaTRdHGqF7dSzR
FIpsErRdXy9fbKl92IyDeoS52A6ahskykzBcxfvpIwPbfX/Y8vxyOKBV2X3RFrWXr3U3o1P9s3mg
3cl/dojOl9PQ2ElNkqFZYzMVvutRgHIr/gdeVSv9U6iQTSl55PsqX6fq9Dy5NBNLL5qExnDcMXkl
Uo/Pkj9IhqFg/2OFPuwAK2oS8umkxawehB9RLfD56SbrnB7VCKt6SW6u5xfoJR/qVTsHLByg02U7
7Qs2g9mTVdjRBEUznAwPd0e6IJ7v02cmua3SkxivJw8Ttw8u6G8Pe1GWYNNDHKRf2JA0yXMGG2RS
2n7u0bTdbdVGcU8pNVtQdGP1fbx9mISEdwi/xOUTqyJoBObpCtkhprI6BbY0SiS43fv7nERwSNiq
jMJMJMGzjDBzOVSDAQ75KM84CzQfLUOXfxoUsSwFfXvTH7gWAnabJlQofte6eBXuvVT0Bo13mvKK
gwaDzs3CKJ71kSAJBysv2OYlhg/6CiPJN/CYuSh0GPgN2iluPuWa4zBpkna2EC9xIVqg9wAXMg9R
Ylu8blwNg6LKxW3pr8B0Ph0beB4v/JOt3tanH0vKASHZg00fe3vFVDDwAQ/mfuWnmoS+9SbJbWWQ
Wx3IYw15k2uQHB/L3SfDJFtYKefFN3L8XtkYc3JZoOKkTmKP2gepCCjr7L1Dyf9FTwY1/P9+PBd+
KJ/77mBIVA/0siD7XhitiQfLDWJFww7zXiweXzDTZgZ36LJNJWC6mI5bebkRX/lFY7Y6CX7URIaW
G2wuB3XD6DUqJRdwE8k4jaC4pdjnNTUiurhkCmQlPo5TGmYkypZVtszPX3sGqffe05Es0Vd5qiQl
JjW2dHJiwjLx6mLCFE/tG0i3nNsWcI8XffdEo2wUVC41d+Cz2T+WH0AdqlXAJK7cjp0y/rXQYXcC
J2Le2tUR+3sRDX4aALHXRXwEeXYWXZlDsRLg/hJfHqodBG+d8uGYZYKERSllrRkj/60LZohcpt0z
c8O9R7yzGU43oQ1I/ZuyjxdlswtTO67nlQf6KEZdsmuayCkH9HMZ5TyeEzPeXWuE4U8ZXysYJWdh
ndfy9tb5A64hEDj6Fy08snpOqAZJdKWo1DGOOQPgqW0eyQBIkLkscnLgGgiwHYq6yLDgjvaArpWB
icTspNwUPb9ibgmbKA8giFZWQiQPeyCITM8zmlJiVmd4/mpRF8hg0PTCjJo0ZXEmyOjsd6lY4XIH
xU8M/NrhLJajRlj3WoG0Pz3L4MLVku77rBZZHM6xHBtJPXBf5LvQI1rRxsV4a+cvAg/ActfhMxVo
p2nrGA+/HK7k1LKAId+jyT37F1nVZOrdHGcZKDAE/67C1zw5C00Eg3PAsyXStVJCY71qW6E9V+7P
npWPM6nu+M6la4wZ/0JV+hA1DKmgplN/yfLjus4JeKxWp884r/f6wnqzdXzdrpSbtN4m292VF670
yM6jEAsAeaBRsCESj32az3Ihr/9IfFADwrJFRQt2qqXhRdF5WK96CJNb1hPI1Z82+k5dlfvDhH4O
WiwO6YstpVFJ7UK+GlB9INMxVQLTTXtmWtiQ/H5SNaudfpTrc8YMkBXWsvwdB2lrpo3j/CzQMmIU
j/bpIgdx2DNEakzusoEMFD6sCTjkIzjO8flm+zVYlByfATlnapLCZOTLrI4O2RFHkSBl4FOu0sME
DKj3Q2Im7w+8oEJAHE1T461VxmcXPZBvfXbr1VEjlOyC9N6S1Qzl2LdeSX2sXbGaNfXX6cx2rLzB
UqJS0Y+SfBRwrkmmQmqJlvGRiJfqsLW4++SdICudIBXoNOYc0h/TJmg8f2owT8zgfmUrzx3SHVlQ
bJu45Ae3btP/nWOQ0ijq+C0mHSNi9fyFFzXFQQnfcDCvxL4j2udBrqT7v8vxMW3xxlwKsJoxaB4U
FFalU2nuoDBjuxPKLARj1SrIbktvOw46RJ6++ADtYHpoPgPeO+gwtfrcnJcno5h6qNYflD/Gqlmt
7fx2q0RX3cvSc/agiRgZlu4PDQzUTxU+mSf8ZlfRNOKx8SdsXF5Wl+UiHKxc/RP3/9fodLyXRk90
8z9WY+Ayf+QJDGuX2NtGPfMwUzTQM2BSAEOSWlNVIb2T7IEGTLHz3DGIjE1kH5ZTvBAr09u5lrXx
BTr2CHfOglyTCeX31aUjlte+9Ig76XqE9sGidD2AWdwoGYlj1Bz4/e4EC9IeTNwIe+g8tmwunUyI
avXlmStkOvPaOLbA7GbTvVfGy8WxMythZjJDGjbVn9HNjsYpCHRgALQ6r61wgrnvtpeYIpLcHSya
bhRHWsSKevfAVCufQpFdfvC9g/HVQ9Tiw/WNIdA3sNBQ3YNA42cjmYHuxaaPlSq65bW0ptEOUbsb
d1kWa57wQ9aidaf2NNhel3OfZZlJ0c63ldOVfZ4o0hM/W4EHkNeKwwmLfelL73lvrb/KmhBTv2Da
cDT2MlvOpfvGF85wCBxBq5h0RDyRN4If9T9iQF1TMd/bswhUH8nzDkNt+XR4O7n1ekyIewNYtnLr
knjQ3R8+UlFuNU3LR0ETHAG8k4okvGTPc6MkIF5l+FFMLeV3IOEvve6Ehd+qhjeDwm5d045RJ4ss
X1s3PFc2ZKMDMjs2BBw3llXFp6/3JGCXS1jxwE8pBkZWLfZFd6Ypdp20z0jaKjYO42mOb0x/+o0+
elyXHctstqnB8JEyxBIfvpMMQ5toSj9LzoGm1zgPCijhBcUNDw2OhlgrJyqd6ENba/qFAYJyS8GG
5+ju8rSOiM3xl/c6Qp64HW+Qw2JC2kbF91lwwWxTzHQuLUpL/hODPiOqUv0aM1mn4CwlUZhCeXFh
Hb6aIpNOFdPG91U9q7XHrattprmyjLI+V1oXzGCqJPNng7S7ZUmi0Gd9G+hNTyRTwH32XjjdEITu
soUP22+FdjknBJklFfQJWQFivNZ5sjzF13uZfS17gSUFbP9evEj0i2pUUnZD/pzWuwPMJVa1p8Qo
0J6Vmk6GIbiGOACb+wGeUEtasBOOWEQpajIKsTHCoKgAYCGYUzLAcYuIssmD6GCUz/pqppLgR9QU
ALcWjYFzFwopleDFI/qjIyCUaLwTYp0qnx23yrU5hG1eHll3hFY+YLJYPpa5EO6ntCu0y5Ufv+Z9
yOabfZv9l/+ewCUvo8KpAjVIi2RdYJ+vImHiO7rYoudjFpk7PAkqtXV7VGb1pwWKPfDZpsEYCznI
l4zDomhH28EK8+keAm7w+xN2I21I4nCucwkI1f7GwxMeHo1tlJqI1EpK+kxyIiTwZ7LlfnsmDpkt
zc6pLPHhZHrRlKUOehSIxXImDuyz3ltvxJPo0X105EMqdWIN6Zcusz2BqSRvLE19RU73xDwnoN1u
Fz8g221B8qKzzbw9mL0GPWsZwAscXR4HmFFpi/HSNsbUA4tyCoofl6rTNJXuZuwbyuMXtL3PkUlF
XXTzmaFd1fM6bYtv3T1qo1Pd9MTUpns7JHuGA94Ukehfo+gX4sDh1ftAIrsqcUwYWqoUW+FKxG2e
DfCYQqshFeFxJ+RUapULpY8cIr6WMkB5m0jSHaiLAj1eZRxr01q3VrLHGqnd1OhSr5KuG/697U3L
0+pwW0Olc8Lx1Wjj2Zw/ehheA8RhNUto8+jSO6mr+JYE4G/KdkzYKo48f8D7UBeKi1sz4utaA0er
ILGDvVVCgKn9+RTqeza9Y6zaocXVBnW4ZoXlQ4/n/dSjZaDp429ENgq3QfTbcRyNOMPr8hmWNraK
sT2i15ywCg+3qwTPAZK7r1x4dT8yaPrim6bb6oJUu6AXccxmM/GVSRx320PZBsy2EKyJSAYyL2wX
wU8CZQ3RjLknt0KIgMj/gfRQ6nyxNB9gSnZNI6LISdTVUL3HOG1xmEA9fqEjB39Bc/kEP/aIyR3u
qwM4fphPBR4Au1/m8RMh9tXFu1HsNYGimYT2aH8A+rcmHF8Mqy+qKcl/rJHa3AdxaPG/4T83AkG1
zz67w8SYuOATo8jja0j/2tZ9F080MBEQEO4dS22lP/YBigt2W1UAQ+yz+JRfRQ1u89wpMBRaEaS4
NMhANRdvcdNKrSP4yQ7xT4GhwYMPaIQtbyW1Kaboq6sThD4pYf80+1u9KO3FwzMv2IQlT34lRjks
jmvn7Ev8QaCDT6SU6exsygD2TWCwwRbZRK+cAB2NxpuP/yT5yIZegtKdpjNvsS4xESURBSHiMwjR
NY1hN+liigtMU6A/+v1VAMs8gXOaBsrqSP58kVsLFKUKBYhA9PBDTOJAW6qQruawLLryEkSxPioc
mtBFzmlARwOf7DpK1iq+ptcpHMVTco0ZTXK3dUAh0QEqRXPxmk3k65imudZLPIjkSSpQL+fzL4UW
dqS0v0Px54cmev3S0ZFWdwUGqbdh2LJq5Rvcc+kCdH/fKvUFuL1vszJlw2xwB44955HI6sIygbI+
UT39w+JgBzCazr2rynwCtBb79VcPbJXHGiUBaFPJc7v5/D61nABSfeUxOAe4ZYizI7NwSaASw6g9
TKdtFSnl0IGDZBr2wsuj55g9xk1oLd01zXnfEpX5FSyBNHdVEZ9c+shy0Fm4wpEuYtnGszglIrVw
vhRI5QvtfqJu49UtD+WCbIzh78z6sWHbc4ic99lCc8TABhA7tqtPsNeqGClu4ggpXmRWpZDkL+S4
3fyS0ObCe2dTU7QziuTv/tya3/VQyhPGuLVi+jg9rU1e1Uzdskbrgu3uKcswNzZMuHVht5PZM6b8
0LFwEDKgsnwKzeL8nD6/Ufmd1A1CZQqZJYjVrdkjQlhb1F4aCau3FC+gGJ8WLeO934bGLoJ3Y/i/
yoCsG5nYaEmSaZgXhPpfrWI2/TpPv/AHumrxEZm1o4npnjNPY2FtJZJYTgC3P9Vq/WXG+Ri4XH05
6+I07UOPi/WRiDdZHHhL+sKosPO8K3BJVByd0Y5OUQ791MT+qNR5MWJzIEum+A1+jepOdOGWp3TA
k8Q0YoTimpef2ZmD/FDKSj8zeylX5u5/Bg0WAtECyP2zUPS0FtN0UB1p0b5Bh6YJN2PkiS9Irwlk
tK6a6uar+eOBrxHBr3lK/5uxH3m7ZU6YgndT1MKkFlkZLRKFC884Mq0n7I7s22wCFMFp+o8NETHU
B/cCEV5W1/pnVizCILOwivsVv7yR600Ig7GIYl8cNVwM+wAWCeDv5OgUCrj7RBCLRGE30iEKXWay
fvStaD9GpGcEhSTLdtjpCz6gieePFPuBumF1imbTmlt1RRZPq3rQ+Hf7FyF/3TIubT5i1v7xmTny
rQSN55ne+cCRR8R29ViRI0tFGIacG9cYDAT+/hji/Ykve+DV66/1tJe91O3k3JhujNxns1kX3fi9
0Pjy9I67pXX7gk9aUdni9MAX3yka1oScoLrcpxNhgZ5VBOj0Pkau9XuWDengg9TvnUcbhM0nFZxM
8pONdcZUz14GnKsXlVyAPFe23Pxm2RmTXwkwKGHIP33ZEScAWIhH425JVWVqs5SxjizSYcfpE/8f
BDS6inpQ+zNgJT0SZFTCADEiM7o4bLPiPRk8GpikSmp62i3wgQjO1BDgPsvNJOQmbgaxwmyeG8gQ
f2GFn6+UFdmPO1ukCE4XLym2wDTkiJu6/nmnsBMzYS3c8hSO8fd9UzNmPn1GytyZ6MMpnwxO+xSX
K+jpG//fKF7/wGnalTZl0+xuOMXc4IVtOCEmj6gsd2wC8RsVY2COQ0LhDuC4kole++7dxow9dUnv
iPeImnNeZi9okArzKfTjdqnH9nTU0FHtJ4zoEiC8Q58BpovbVTgpUruR3WIzOFJTYkgoJn7RGkg7
g7xDNMlxFrfi3oneT/1E6q0VqsoncT8v9OacS6H8NtHRwhmyWY5u9gEvFf1sV4Xi019bnqome/ZB
3HFTThbgQcy+r5srz1D3qb+ZfSvLqRwItsrhIl6lnxEFJZ+cmQCixSZ3YMofl/PqoPNQDXVIpxfk
qxX/EinUUPziB+RzmozsHjtF8H7P1jUKFjQyYGG+3KbcrKU7NjM4eWAbOEZBN8VMuKVrqfgLyN8d
wc2Yjzu8fGol1CeDPqsywciC6oWl1WSqhvREmvIz5C9hxsHViXwWv2Z7YRw/LF/449GuSIllcee5
Oq+xGqtxIeKli2qgdexchB6h+AGaZaA/+TNL72bz3ZMfgVd1ePhuoksD9AuuEDg96UFYSV4RPJDG
Q82FLJfxu4N1HqIFY+7i/0rz+6fKYZHkgsyBIA3NrqhzXfI5cBXV5d/Biw/uUVHqrbOoceXTVvfb
R6STU6ZAjJ6ejhHX9mYqNQScfhTJ2DisvCbYc3eE0vW1M7vcqUH57g4uQ4VB44naTP7/VeHa6yRD
sEUDJh0KEwalHQ70DfTKPIP5CWIH8h6ZEVgb9S0BZlN6XLbeP0+g5SDN7hqtU5csE5/a4Z9u5Wr2
9r9oO2TbVMWxwHY33HN7lwTRdtz7EBogZcUoSpjIgFKkfR1hd9sHLn0wvMe1oxpw2RRN9APItptn
3SfxzqeT9smMtV0h2KPP10oV5+XWePaxNVlnfKeVY+eaHi0AFc3cPSO9jamwKJTgqkAVN1jhc2Pv
FTAvPo1DTr84YAxa3ieBKqInIH+JGjfGH4/0pfSeyeDfRXnH9U86GaUikRtADf5zUg/kQw/afKAl
S0/AMtQndhfHqf/HwM8zRTDfjrJp2I8DEeh9eswJUmRA6JEIdK4hQuSuPP/769xbJQMeUymUFyUj
xbE5JzJMSUC/JJa8bdKA0bYsey45Eq5mvh06Tu5w4ITdtB8J+4bXJvmLsMWpmVl+ZINtUZOJPTIe
DIFPVj3Hb0DKkpHmPlwxp296Gz/yHnDzUaDtoRTApSR6dPiybs1MIkel5MHUW4MRTYOer4NX8OUQ
aCo9rlek1mu/ysns3/ZFaGph+eiw56VuPom3Ij1V6tAU2jHxUvZ/5uCyy5Qx36cVaVo0X1t4dGlN
JQJWovXf2jK8mcNcLF2VIAahTpHr9MsVkDDEIgzALPANpE4ZM9tBtXHyw20sC8BRZYDyDKadJD6r
5ZPtN22BqvcbgsGXiMAxzaa92lI1gQ9kJaRnKqKcignsfoXjVgOzQn3+1R5sTl+qA364snnklfZm
jLSvlgO4feCE+eqM2vfnM/DG9tNBG5t8AgWIRz6CUn9CQ4pTHCclI3X7wY6X6iqT7ydBVr7qLX5a
BB42VmhOjBo2L39izE6Ng/86QBYqFiuKuIyhnGKlx+JTu8MM7hb3XV/JXEK8jlCkP+dPKP8j9Qqj
BIXImdagD7tH7vg05QfROGZ3ixiC8ffHAlHDl3HXDqjWU2yi6ho11PINtXvThot/cTOmyLAltlX8
vkssIXy1beqltXSggyoT3oo0ujSnka2lYcSAzKzoHUOEO5LQ6ueMns+QZxnvwfUnTiALKaQBwQ8A
Q5WWDwTJLW/CVL6jT6hafJ9pC2tkGFv7PaCYETGvth6AvGicbO062lQerw5JRyC4pz31c9oRpJ28
IYahd5V+LWxNRr5Su2Xu5qEXs75HwSnLbBjoL5EKsRpvbO7MgzIopzcXbLxHuLEGxYnXroGwIt14
4dH2Rp4aN9STkwbiK9GJ6rpwWCl1jM9BQGFXlg2Nj+jmjmqJykTsF1W5EeBHCzMmi9IKcGqn7xCQ
LYoJJ3xfXFo3MF/uOaBxq8rfxtoWzl1EnAqYpWmsaqcYfvXp+xKVFERSlu9hCRKX/BSy8fx6n+XA
2IWP9l2jvoeFttBzL2r1DqIokQ0t7UpwRxVAIbq8+EsaDxFeIAG4k8ZAZ+/Qjr8d7FUqE3VESYNX
s1f4x1iTG7vuoHNsvkBAbUHNg7ndIBZ7NlorhXz5L14f3WdWOzC4Pfty3c/LAml3xQnTL9f6L3Kf
3CtHFv2FrXxEC33jW5J+n+TzKuPsdUYK0dgWuYJKbKzPA3trRDe1YKg37/i/hb0O6gDjzHTiQ6or
wfVu9Y88XMad324R2yGZnz+kg5h1u+j5ZtbpL+rnLjyrB5V/GQChdhpnSXt0AWxF1A/S3RwG3Grn
iNBFtYS+Jrsdg2G1BYQxEYejgH6+rLr4JU6jI6ql7km01yP1y73RM5j8eeQEY0ldqdWEha3VJCnL
2t7Qaf40y8kTjj+hM0E+nuW9LT0k9W9IjEoIz1DsSe0RCeRalmv9QSz23PMZZlre0gzYgioye7fh
hV9XIpULSOJ/RhPufvbH/65ovqLEItJMPv4O9Orsj5ksWgve7YVQx2SYwoATwctn0actc9Z8TqXR
1ntIWNcdEY2OZJOg7jFmMgsd6tnt1jlXr8qwAcRHIGdGy1xlYJ4o7NnEquEpbActNUKL0Oisma1R
jxosgHMtW9IdNCmGylR9Ao1/HTPyVj8bHVUzNt+nUfy19u2WphJV00KKILt5FNH8YDwSinKnkl3P
RY37z0dAWmh0kxwCPnRCbNUm3db3FfelhQwoXTMgE95w3oftawZ9PFqyxrxYjOIiWA54xDOd6GNB
+P7WKsikSsQpI9s/ShfNePYUx2YU6Mf/wfHNcZdeoltKW7rSqundSjsyBO3vptNMDhbu0e7fjxD1
bRHqUpfXKaXy/cIppdlsM4DL4fEsfmbgYayyO00dZ5FsBMfMZjcczXBM352kNCcu6UkXJA8Yf3C7
AT0POc9Aw6FHhmFYfT7Gm6LDuKtWot4vHLcYmYeQ7A6rspaMDnbQoAqgQTuAJS/yVmv58VpHW992
MOcSOK/Nibe61kW30oSjuDasWhQSQnIwvsPiZ9/VU/oLjAC6QCd9AsGjvigALFNPCzfTIbA26+Qq
dWwpBNrYrK9u3qE81GGUj1Aqoltk3dv9oaPBUW0KX1AP1w4gWV7o1PUnDKtspEv+nUbq/HiaNalX
qArpzY6xaKLcJIK6cTOVWwYxUipgVEeo/sYDzF4pezQMZs4VqP9/MAa/h8/7QjADxJIlGC8jN2pX
SJWZnJEnThvDf3tJzFMnHv0ebA9jbcevr8CFXLaDCUy9tUWBC6ZLUtKv0NtWB+w7YCIXp8oVzpx2
QmBmIECRBmsBTsN0k5WF081Cb2uZlIuOARTgYFuCZqYDH8zXS4jJrvKvzfiTgjKOUrDqfTo0Tpgg
KVZsXt02ia7XdJwVjME0SIVc5i7/XWhCNcv9j9wnbY3K2jRGIy5N8dPgDv6p6wM6SXicZGK5GL39
vAEbXjjSden9TOhfJFdGt/h/kLDt9vf6O5wJMAElLjhiR/Yu9Q2dZxTkSGAHB9zUwGcPud78NJ0l
SqopQ55PopOTsFegX/19EqxlZEYHTphZDVcd74m6ln1hgpKATX5JRX2WJB3akfu+kW5Hp7Eptynh
nf6rn+zzIffksePkXSWU1LlRWsGpO6UM4zwcEa+2GM2ckF6PQSXDPUMkQBMWAGCkMdVYS20HOrEB
h2C4UDERnW/3Kljdjc4A0T3NEtxFQNVCRy+ze7oTTLwUxh3pEGEJjHszVMh7Y91ZqIpjKV3cuE+l
ViFu1ElVXv2h7hdHymVDOavF9DLzkMUwJ6XlzlbAiDtI8guWQjCdNHxsfJeyhVZEsLct5PfBDcvo
sVddlWoDh3B1Bju31m36R6KM5h/ieGPemSpDw6hzUnoeY5h9q+Df33PtNx0vleClIDtkNVFL5vGQ
jIHvI1a1RTs9TQg7kSmj7qNr1d4ookNW+fPFbtdtBWwzq/G4F2IHf1JhHGKnpqVGLwta5TarX/7n
NhEgAiPvobmLU9sGVJZmVKTpQ2EaMfP5aVFQ7eDE3KKY9R5dE63hDfC4YK/Nn8modSH/0MPYickI
2c93Ka+nYGEp9RlyUPC44MhSZ5HtPVV5LZJ/xFJEv+cItK2BmB2KXBSTGk1YgbihHly5rJP+/FK/
Q5xBYs30JWjG1DikI4H0HQvY7IKvvP4sZWTgEomMavYgZdqqzSgbD5tCNI5oOMpMmt5FjDqWj4cc
NlvgdXWLbYXQ+ugFeVe5JEKaMV+RdG88aA8eeSAzRvwdSkvH0NgQVlsk1nAegA2xJgX8t+N4lWRY
FJXNIg3Kl5/GSZEe302xpND6EQym+aON1bcLZ5IWH6wcthz2R1Mxy7UG0DkeiBDoWbQtvC5D6aor
KSKM+nLhQGOHrmkx8I4cUD643nBQ71L44Og8JaDWVrq6b3Ed2f9/bdL99Qs4R0bDYZ1uOa0k6kpg
hbaVG3J2AWE66DoMgqe4yM9A09sRjJ5KCzoQmQ476H/ziCLJYqrAWi5H5xQNRAC+vPXmi2HHC8Ov
9FdbvPn2wi7txgkuHpT6IxavKXhXzfGqRigPzLq8lEt8FK9Fp42j17vaBZbaoWqSiRSHxKkbY+O1
6FymOmFgL1rDlJHqqqYrbzeXujiZEekuKOSZQGOCZrXelQfCmP6k2d818uJaVlqHTiEu7lxYyI55
KndMF/acb69njkWLamPRKW1aj+vE1RxuJrlWrM5JqiUHiU/e3rI0sgeH8xmQ8rwoUdHwsmACEUp7
HRTE2ec+h1cx1k1g2a3ZzkUQs0gLnb+xMU9WCTCqtmTXIhgKZ0tK4o/ZZvAxLadWG/BSyFrFz4vI
dDRW+iuhkIB9QCY8aZNi93yuy4T7dYRLvHEdVNwdqmXE79g0ZGsjEvFD3BVzjyQ1/dzS50AZO1xp
v8PEqLL2NnH03xUiCuUghn+oM3wHNlE6CWESryn1KYL63Ihnh8joJ5plH9Xy4ugoLQArKYPX8FVB
uGiDevSuwpagKrH6Mq0IhxqM1jlxY8/naM/Y6rZoaz0VLoghVccPj+ohRwYrq9l715094BB25PLD
ViHBY5Wmpdwege7cJ5BKoCSicMpnsZDHVoroU/5ymAsqU9ZMgElHnSDYcvUxXnvNeDRTF09gm5/F
MByNdlvZRQ++4DSmfCUzov8jR6KjbpkqLCJ6Erwgr0AJ3hEPmnx1O0eZ+VvF2oY+LurCmD+PjZy/
w1ETr33dZj8WTMBgTVhJ46xf8xgfADfwXrsvJeVN4/92BG5pNW8fhcIGV2p9tSScWhAXOoDoxGwZ
xPKsgWvFDiC+StQjIZeWWb04s8cHbWbJX4aJRik8AyLFZgYZRKHXpKBHAmSgBecAadC1bBe5dB5w
LNjrIWykJgIyxFHx8j3GRdKBrXGpKjGPBviMuUt3PveTSE0Hv7g6/vOYQrvGwZ/COvAGIMIN85im
SAZWTQLkGrgLyPeRzO1Bcc+ojq5QfmP6IqChOcZd4T9MqsSswDY+aIPj9sGyrmiHqVSYDeuV0KXA
9EtZT6Q5XxpVseKdFLrEFkgWDoqCEdZTzTBl0k96Rdn5s+2to8HzNSYSn4073seZLlkEWJfMyyxP
Yzc3XLLVzm91XK+YLPK2zbg4ln2iCQ85rRJLUKLfxYRkLgdqQ3suZT8GBWBbP69mdFvrb/+sYrHP
AeDypO64rbbTZl/77Zqwp1X645iJh+7P2ZEU1W3nXqMO1ia84fWmRDIXxOrh72gq1/7i7owvNII/
jGzFulOgO1hGZY4iNeMWOCekcoXseyaq+MiM/WwfjzynYso6m+ka4SDA4eiCmModsWC6K88c9clS
5LB0BcVDPl24PfgjOqHMzF6UlJPSFNPLJSYe+3EtAgded/YEUznDNxSLbR7mXu6b5g6OwmX/dTYv
f37/mj6/c99nIg9T6lCbF5qqpfBlBvXcOylyGV9oMz2TXGYoZViTtYoi/8qQwBt9reW+/drY572T
Vchhe/MbiQdnjVgzjrl/Tre+CwS0/Y/fa/FWnrHH321Y1uAwHhP4nV0AcYq1Lnx0iRG3/YZYhu9i
cGXAqXiw9tILlNWaYHtjNSoZdGeCME5db6+xQ7/shZ0tySCa8AspQkqD+UFvMLHRzku2IiZeNC3Y
gRSJHtLvr/Bnei3ostcxqVauDlbLHTM52Ssc0yaGGr+e4LQJfnQSIjcJdnRP7cQgsg7KzIanhWRz
i9u2WwdXkapKUpaewuEwbd1gWp1qQUAQefNBo/alVlm+w/HlMxpF4fVui2Fi3OkxUD50OPIW5TIt
wBfzaKk6FzUnpy7/9MYPC6V7F86g/OYl5X7KLfEYXUqLnnkFVZfy0xv3W+QE/glCGQUPgXVU6s4n
Cg1DY4tPsrGRq1iD966HiU1hILNqL9F/GICYRFGp+Habhps+wvNW1yprE758ssxOC+SvKjcx7m9B
vUjwHih19GL7+YK+lWBlqoGu0R8miaPxXt/JlbwPnWlRewZxJ16Vp4DEp0cX7Ot8jetWoTyA4D4N
4sIY1UnUaROm5XC9qCZFcyR635MvNxxu0lVWTbsZjwGwB4xYOMkwvf8X4KGHmKQbXdFDqH8p1LTK
1r5Dn17rBwXWXngZTHZ25pWrZa/FGxdjVQ3SKy9lDMYJ0lw0oeHZX4sGCULB10fUARSUNeyW/e3b
hfUBc7iWcp60ohOSJhBf9NyWy66KxIZuF4RHiXUijVxjy+U++eKCDR/oS9NnVSdhmy6aZ2czPrD9
JZvfo5qXWTZLiSTapGv1c6yiMY77PdUVqc11hG75x+CxUHZ05KUDXWkN9CuEhxL7EOarHkHY51mw
PaoPt8mGdrlW3rSEGDZhmkNuiWQQWx0gnUhGmmleUWeW5QLt+4+D2cL21r6fv+/6S55k28RCLCLW
hpPHhGn0wFCtry6k2XgYfM6pInEE9xIDNeH5HduPJfVkHXRyzQZNZkFtIzcNQhf1ZlcevrbBo4ho
uteaUPO//qqMkWHY0NPo11IltoeOooXM47OUXq3zHt7PDkieqR5vTfi9oxXqU8JGXhedqERjgjfJ
BGrlze+lr3fODeZikddwD0IxI8Qb00nkSI7PwSg9rBBnfyM5GousSjLCRstOn29D4YPPYjMzRwQ7
Nj3FGtSDVAy4kzv3/SQbi+T7QzwXYWqhFABxAJOeG1zGxBvhVzUQ5wV+bTw1gMlreAIEyaXFrcuY
qjFslYM3tDRMZ2T1SqXcdUQIi7euT+xqP0Vsqui2mOIy6gaKc0jK3zbUi2xRfcYISYAvOvqP8Cut
CYfeAjE2b/Q141kXKvvzk/miWvqj5zi6gIILM248MCoeLMKePYxKlED/wmZPu5YYIWTIr0B+uJ9+
rHsjmCPv6m/4mbmBzXqrYnqZFB7yd6i1TAvQN27M8NrdeX9LddGTG6+kTjQITSr74E2zq7lw6rQr
WOy2N00BcUUodCIjWnT9+WHsaDe85X/triNZkSivJKEIqty5cr3UovBV874mymHgAB0WGXnmKtw1
CCgz+WUAnbk7iydacfd6jgbIUyFmisMXzg1cimrDeAUg8MC6JYoVH68bgZqRSlgiyPTD43sbjxOp
05AVkQy9ZJU7ZFcpR+mdArQ1Q4vJYFJwglCnZ+hpnwWsk78d8uRgn6KVZJSGtPYKYDiWHoAalmpu
rDpwRzcZ7bYliPCN0AiGvmwzknjxw6rgcpq/xKQ0/8xxSkkZB2SUQh/LRs8JRCIXziKS0vx/0bSg
TBRYDWmwRU/IDosdc7fZNy06L8ir/zsMMGPeP4xGRBrgxDSM0B1dc2KiCWTag2iuguaJ+al0C/ok
lX1cwN96Hjg5+Efae+t8+gwhLSzm+X3D+8EP8U34fXb6YH57XdVZHrNsW5fb7sAxODnGbde4zx+X
+/slda6jUn1+lvLQO5qbVzLAUlRkoMLuRnBP/tCccDWAzqTXSG9ALMmXK7ETliK0FNx9wVt7ECf1
PZwtjYkZ4k76xOCJg0fBx4Z2JR8pbdVv0L3cMQz7C94wIl16+vniJeL0iri3f0GWYjV88mGIyjXL
8eEUS3eTDWNWEufJXt9WyI3VtNQyrYSRBUgfY44UVJa7LnruULbyV7u8BWJfih09tyoHd4stzfzU
dgHbHqAzKpWz9zUmF1oIWcBcX0xmEuzNGjDGrYa38xdFY6D7TvyqFgLB3yV5P7vi7oZIdcKWIEFC
6QsnQWjOnHTAn0eWh786tylN/u5v5sMF3Tk56wThIo1vUpqKy1UQDvWv4I+nV/W4t+Gs6DAVzGUG
lYnbWx7MQc6dIpQYyrMPCJXkuzZ4HmvM/mzJNDYpLKhFVkBCQj2baV1fb6doaL7oscyhru/o8/OM
QZ4nUV9eow0kRp3lwUe6InimcWNkgq9CuKnwZUo0F5bbgFf331j/UjHnHLYYv9JjbL2AevLSThzm
D89qaXAQ21OYSTw917Jl2Ys1RBXeh8r9pROf3Ch6Vqcb1BRSo8lwrOSv3JoxADV2LAvT+t4INjQe
DI6b+J75x+RhVB98sQ89B0ddiq6Za8qAwmILjSjrrUgoFfWErxkJ1p3ldxbmM6gwpz7SRiu6jQl2
Onn++T34Upg/NwTUDt9eCunohRdgpY9eccG2uL0RmFtHu4yu/rINLDg3+dKHM1BYVMiR4geD3F9f
Uan5zl9uVLpEnAMYNKK86mLrGdIZAZIyq5RClJApP7xZqRk/DpNW6KA9bx1ClKNTXcnQdL2DBlZN
VCs8Qiyum5RxSDbz1xH6y95NugKAAII5q70+mm9H9+7pY59QstXbWMyD6xglK8IQ9tmZsjysx9OQ
WNPQkmd/s8S+NBHyMjLUn9FupcbFWGrgfIgmbC9G6G4GRFRkmVuaNROEEBckXNJxk/aLIljcOpTp
Q0pJ8TH8jAOvuNhr6fnid24JO3BtORAVbAo59hWmIwgRlg2Tl6ubT+jiPP2SFnR3xW4O7QckWZNy
e9C+7ijKVzK7/vnGJszAGt70i2LjMHzwTfGTiuh53HBvNKf1/uc2+KlQFtlABbibGzHyEaBmJ6u7
gEgbyjsWPhjg0N3qHcjUG4AjUEWFyrkDyn3GlfyKuczJ6gIM4g194WQErEXhnuJD7Ko0NuAut3+y
NaJig9IexYxdJb/Fck6EwPLSQ4hgIDRZ8UwX7YmWQve5iqyfwx7GpSuKwvazyK9fuYIs2jRQJQ5L
yux6gS9j5xg6Jnc9cl27YBCoUNAF7fHj0Kqj3pVLMAWjM6YyBi0XZ7tRl+lR5+VAC+noOH9z6/ld
uZmx5JIruvDRMV5gfKHCzz82dAm5XyWmK7Tr5OJxqAT6cXvI+Tx5tbp1c2eIaY8o4heMXZ4F6UMx
RXFdoo2Wai0M/iBp2OlxJsTjhw+1Say5BoL0DHzfnUyoKSzMYLmhWk/N0dJq+QSTU4h+8ENcw4O1
dQYYtaE3mMzQcS5RtKBqRX+Lg18h+XO1K7OAdxGZsY3nNXxY8Gj6O1iG5euxpA4XmQ0UWJ7oJkZv
cBNCEIvHRoAL/McYAVTT35ntnFARTt8VCyb/KSfgt6F36K0U3JSQDDHc1KsIh8DjpNEwBBNs2bMr
dnHJ0kr51JCr+mwi/DuVKr7NWQuAKBXRUYkyXVCVXuOvqeOQ1Bo+Fgb/HVxl3jRc81XrVbhMP8s8
aDAWzXYni3jnsgY3lNKGDcTLkOIDvI23daH36kb/EurIKNsYKy6qXaSvakUMJw6XBK/qEi6fsprR
xsp7V2J0TvfbkDKndgKuJZPGVW3biiW+kefAt3v585OQeIwhZ8rO12gkltLnU4/tkqevmV1VpGv5
mF/cwYWTbFGSKbyAFdwJ8WSnQoZM6QT4+imypPnosQssueLahEM9zZaEKeCO61Tu9dXjdxPyFCMl
qoMIcyK/9tXfaOrO9VQF6mbjFpwyz+tD4+OtJUzlGaSuxzp0FgqlecXenEnaXC2u+6+IACLA+37t
TdXqD1knA1FRIlIOrI2kM0GtSedaz3McJ4PwuVpegLUwpWh2PWDRQ9tpG15DtMyC3J98nP3ozbSn
UlQXNGTM6BV7bWh2SUPeGQWqWHBdTYQyQlXqTVsR2hxQMwnX9RmpJzJzuA3QjC1b8lLuws0rTJcU
eX10ZVsqagc7mgZNpwN3hNYhCBvpVwQmV0NLlvpWg++oYFGMBaQu5xL7lc8Am291NyeXExJ4F4Du
gMqwGcR64aM/m0cIhnby2yAIA1YzznxdeYG8cJGg7q4DXFtvRZl5JDjgnO/bSe29HtGLe0ofMa7e
BAqS1QEEyfBALeppHuFbJEnfKywD8u+BV4pTZsjNjfFGclFwnkqPWAipyUMyXvPrTlBWH2NhQuTt
yXMGWRt+0kUmKOhEKR9dCCXHBZBhhf6MgvhQSDwl9BYMJyTibPL+faxs850UBOTFQ89axKblSXXY
JLFFmcydC4XUZuTNHIwnruSh/re4dB9y2InyMQYRIN5mSjZ+OiMgaFK8vn2g3gcWbtq8lzqwbARf
H0tlq86/m1BGzZSbehxlmc+ZPYMxE9lRaNBo2SJx/ihsMEzPQKZWPeJ8z4lMsb0UkGXdKnA0U9EO
1ocgM2sbhPAWgyKLffF6S0rGV+MysbFvhWOWNfQ7ePXkAztrIDoNP46+C4YL+bZG50gVS0YoaiSk
+ohr0wT4odhNu3blI7VklD4SvshZ3fPuoaZfopzPpJPl04Tb8OOMMtjPMHQ4+3NxnGNAkLXgZUZU
3xpDq2rGFZ41btohQU77glU2t6Ycy7iy9j5tAwdJSkCIInNV4/2cSf5zYNCt3eJfndhAZpp49zn+
VLv02eC4nj+D+slEeAP8HewQ0dSN99jSsSnmmvZbqlhC1CJqEkgDvoiUYAW32tlGD9u0pw4sJqwE
0JxHAGzeDty7DMLHGVS+kf+sQ5POH++SYzMFPs3xG1o6dfl+HGwtUBvC410iPqIG8W2VihuySBVR
eZXs/gwNfQwJ/+iWf3CzlRXxRff0SlcjDC+93q1GmKkWCVWx8c0aCdcZvOEx2iAfcI9FIxdwXQ7o
FGqHLKQdYxG4z8H3vCW49oc6fSeGLwx3YNIHa5dWleJe2z7kTW233Ti6GENaeq4dObYQQgAhimom
Yb3Fyhv1VV9aZCOXiGjJm5JRCHuQiZY8xH46xnVq/YoL7pBvNliSiUXOKQPQ54t0vv3pt0QVgiWo
mGcdIg3vV/Tr/NBS048EJw8BLS+Kr5kWO/JbquEeS2IlpkKcgTlLlNOumVveEr1ZYmpxvauqWBl2
iMDC5pWKSPpKcsT+CunUSjjUiF/U9n+5bkTd2xJ84W0dxsReoS2Ci23/cutleiOppp4tLljkEGlZ
HBzcjMQP6wibpVucfO08Kek9kXGWMxiMEjjQ5MCQ3Brgz4m7y6WSNDuVfygQNhhnjk5YStRDaGSP
bYhv/pp+985R6RBGOnMxWj2PScCdx7GoXnXFUR9EK8Nx81o1TgM/UEOidDoqWcd8w5OiZCDHrGEP
w4GFGHUeDs7Ii3uxMLj2PE+UzoqKd3pTROcUCzVy6hAGNF1UbaFVt+FULtHBkB8I/2e3AHYi99xK
tlg75qz8wJ6lzP79xXZriKk5bI5V5WS6UtOt+rrQM3xxb0X6pZB7VBNsMQoab0QMrPJPF/Pk4pZJ
FL90Y6b3Z35HYYApdW33KQxdHD5WgepoVPG7/MSyjFI7B6D8fpnrwncN6clg6iOm3ALLRSru7bz4
Nay6yJVTNUcp/akEU5XiakwyOCwfWdt5P9msVtKuUjR7ZoZndPRge9uKVchXXyAZXDJMjWHE6Iof
wKnp9WXVwyzkUxDVMzKfVJp4bj5iTMOFP8kNHH6Lo+KHmMq8/wBV1czMffw2e3oZz7wfDesBsuUw
CCvEPuOwj6Yl1DU3D8skcTcUlIFBcyxre0iY0XKd+KsC3jX/7iW8PDxn9ZzG+4e+OAlUEMRjPrdk
WrxcxVw0oe9VkOZ9JQUh4czNEJ7FrzTXBooBKHDEFNsUbcj/396lXk8oGZq2Nri0iwKsxToOXYiX
Lw+FfdVqrn/teK0uAoDf0XPzZIAsh/wxRsynbe6EX8Ydi5GGRBWYG5bWYdlw5O9gcrd06XuKv8hL
fDMokrc3oi/Ix/Vf0T0hkpTluQVD+Ry9BEfs+5DkmnFH4LFy8c7KS+JsqiZt/DNZqdHFH2Bgh+3q
71S70G67fYSeIzGe/dXYs6n7fypG5qXUOaVpJPequkLn1hmim5NVH/2YTixFn04MZOW0xxIBVkFl
IMzboiuhB0NIrVu/hJKxUjMCvyu+IRYWA+D3wMs6w2jzq/y7Zo5mn1PN+06HIsaqOuTeKkj6xSnK
PwKwrq+RXJX/dRwlN2nTUxedC9JeWPdkwqIvq14BdAtvzQDjjSb3ivETEijIVsLWRnX2TYc7XJW8
8wwItetTHLVqA3ZDBjqSo3GubtmZxB9JzggIeVkJCmy74RiL+U+1yt1XQPzh5KzJ69Js45xfD1LT
Xeb1qBtbmHMiQOCvu4AOl7i4W79G7PRgfEMGmRiI2cLfSzY5dUvXlcVxATn1q1fysG9hnQjvyQH8
QT1oSRt2xUQnZbg3BD/cb4EfTxYc7z9+T7cLcPhU4zStTnfAnzgZUjpHlEdcazQP5oN8ZI7+Vuiy
WI7Z7Nr6VV58NLWajQvKJjgqL0IT5d4j74t9UPRFyz+Rm2PAqnC9az6tg1GhUUVIBMT/OO3ktRpN
9+uxebTONhdDi3Q/qf0nH8rdT/N214q1B9MtZT3I6fPQ2lI2OppJ96SEfN0Snhgty5oPvPvhC4Oo
k/gLmLrB61e0Wq/OUYwLIPSScUC66SjVHjKuywG1/YlVQm9+Eq+4w+EslRFYlam4+Pavd0vqF5Nw
OG73SBVc14AYU4vMzan8CKF3FGfl0txPaxSnFXQyhtlXrHVnK1Hlsl5LdCvbt+pwGHc3Mtu2XLSo
cDbGNg0WdySCUGexr1BF6cdir+No9Bjw60CpwAM9Mt0q3lk514nI1vAfw1Kc4lH1p/BQtC7W4a8u
k+/FT+ywcv3afQA/7eQnLz/Qvdrii2c4O6Fl2OcZlvVYeUvZaZzRb8iZ72PQ2JHtDhY3ab1lGTfe
y6OOPBif6lGBYXFZxRtPFQFc0SyCsZSAI0a9GcOhsTD8LMvnd/dJGed5BBPVfx4Ctq6vaapkiXCu
NZFsUfs9NHfAdttQOynZkadDJlq5mRGejY54Rw7DHmYiBPkjSq/dvsZS0xnU6tB3XdhvlOfCVao9
IH2RNKE25ymH1zLiOFLgvkSD4Vn/BPrrYo419apudzqePe34bixfuiGlK1rKl+W4r2jbtmIR2kTU
Cv+HYgXtqYyZkS85H3kn80onoDu08CNQXioRtTsrv0PAukA0j8z0eAdHPXiHbAggojwFexR2VD32
SSM745wq6SvtCorBhH9unWhQc2gvCSa9XjqAA+RVvcmdr3VShhiApFqkDzrzRTBM9s/gFWZSj9z7
DqwVymQ96A7ogc3IpC+DzCjIbf7iIBqzj34K7WQc5JhtFLroZRuVpNOmK+S8l1aRU9rCi3yjdlJW
HMsoO6tAb2EWOREJwmwsp5fdlDvpj8ktw8JfLcvnx3lhCrnEo8SBQfUg90vAk5mi43+xbd8IG4VE
tfskXbnN4mpMFpdURHkaoMEPKVPUardYmBIG4vtTP9ZltsCQXJq0kP0vt9I0+DTJOoSbAsxBaj4h
DtQI2RDgHLHsL56sCrGbTD04k9a7tp2jOARJFn0GpwgpAk0bMpcoK0jCgbRJG66HnU9NS6Y0nwRZ
5o97N0FYjnzO6krJ9b9Up8/ZNfnEAhCZWHwOS2K5QEpnZjP+t4Qk2HxPS4GkFGvXqyqqOWeql1IG
TagUtV9I2Kw7VPWo34qFx7/QqlnMb1yVcAWWi8RqcQZ5EQQ8LlwLfiNEZk/K1++nemaCBdDP3/DE
soFMe9CFCYFYUBLS1IJQbMHayo4Tg4mRJAMEtkhwBGSR9zZ2ZtTImjR9ngSqNz7sOZFXr38hM7cT
xFeNno1SXPYmuZs3YQBylngiPAVXHjLfVcogiJnHvtG+3AT4H0QBqtgGFLZ+K6ZfwyrGoHcjCYzC
OXopbuwZklkxAIauUUFJXzzqrw9lKSuyTRYQ6gVaD5U+hcFpOJK9FWjiqSo+7yPfgKSYYJffqHRd
0vZaK6/tcrSkSRS9GTt9fNwQtHTNPtOmxHXXQKjp4cxYpJPqudEFSPc1oQTEUgYYf9tYH+hBrhNk
S38IbtwSfAplgndXaw25up1889QsICOOEgsypf7wJ9Rggw2NeZpIvL6MkrBd9Z+nXvu29r2tg8bD
nZ0ohnh4/cdTmvowNqSLlTur1jz0xEhoUhjuL5IVEHea3Z0VoLzl7to8vd4jVEDru9/meFfvaopC
oMAVQbKOiSy4xcTs5TW1T05JUvh65lMqd7sU/2LBEz8Z5RzlrNLewST4peLUflIUzpwHhGhtYCOI
Qt0XjqDxRH1zXnTBdDu/AgzdRRPNiyOKfrFeZ7Npaf3UPdKvfVFXcIZEY7KQBIrXiG5L8QhcAbXd
sa3ji+2b6VaL88V+TZ0Unbvbt9CSu5FQLdA6Wem9GDVIxtOv3XT3AfFzOihmdIJxvAPAR04Nm+4O
PBLn2M673JB4dNkZ1PK7O43c2xKXQ5esIiynhUvnnN4kGmJNLRGOQvnTb3UxLWVWUD34g3g6Bqjs
alyQM10kJqDlzrOjQTsHMrzvIZJ3M8f3aVNSobp2Y7eC85sLiSJaYddtulEkthBk1zJKJdHSiWRF
GOzUk/xuCNzHt03CLhp+FxImLHiuzxEZxgGISRHwUHwDCb09RpjTyZbOyrcDGzFILEFk02H4MPmq
xdBDWcHXR1aM1MfNiOCx48t3gjOclmVRx5r0ei6pwQPM9DlhSIJGttX1jcbRY92df2ycsxloP3MK
4/yB09aFT1MMM0ePeGsiBP+HeMGE6etdgF6subPawo8H9y7sEZJfZ0aLvZOydkFNQUA0G8XcayBU
BpeCaisz5q9CIT9fhNnivIMmg0hXNbpFT8rn108uGu1GD05LO8q4gajBEkBgOseGeZzKHIwBJDTJ
wDnpidCdw67ggzqq5V5rtO4a6y6xcwCCO0hAlgGwh5k80lRHQehtHGpXiUP2cCeyu/oLkDiquJzb
jeyAhGmKyQsvRBV857WQfPOfumEbhJz19cF83W4kn1mNPaq897gIYiFSfXWqF8Nvp4PixrtuF4/b
Y1lVVq9jNzliaWpKGVC9RJJEhuQ/hnCh7insmjyUGxsZnQh7XJypnePvqwrGMtq3guMapphtJQPr
85aYKkSTBHX/Hm89R2OqlBhBsGdev/tfoJ07HILE29MnXM2T0Tm7fboyLt9W+8DSoAVIR3bjybeO
Ml8MSBFVjF31EtGEPMATQsFMLdRln0dBlYhLYqjGBviRa6oAo9YckFDUkVcLuei282C8B2LslSw1
0uw2MtM5rnWJQrWZlq4M/JhBJfh3DvG8VWEwJ/wZjE7lv1lwaH7j07gZVRHyrCrON1ZC2X/MvfLl
3/A8NhyNZ09XB3nWb6hHLellcIqcLsqE2N3JU6AjcEyX14mzO8LzmwSxp7WSYnauRqknmH7ehIOC
1xKEJ8W8tkkBevhERw4FyCfE2yBL6ySb+5GhCdcHM+/ZV86wV5jrS/M44vFMpY2wFAIaEu5bzSo7
gn+lqhBJ0ATCskGUWMRTkhKU0ftsshhHSl+0n9D0GZ+ZGmEsBtxqtCLVQyhgiyPYwWAvwUgy5T88
bQ1uUFy/PcEYtpNHPbvi9Fetn3+OGhcOtm//vyCdKv5vHBoUy1JPgzwniyF0nyCGYD6+Wu1z5Fxd
KiMO8kLS5mq16hMIAjhXV80HQlTxoWybBjUkKB93TrUI0xIvUI89hhRMZR4hhW7gF97dg1HMAZdy
ZhQOXvAbFkGguyZ01Jkn9gEQ1Py05MzDrCaoUXSSu+Ie48tK0VPVao0wrHyKM+C+rn3qaMgZi25u
fH6m+hqSPT3u0GWrOhRjtaSkxMHX2XEi1HHm9dFVYVGhNLOvbuGchXvyeoVaoXsbSAZLYNk3dJ9X
/vvfvct/0bGC0pDBgkHqrBlgFPQxTyzJ994SqDzQKkCIB37i/h7BY9dVYAyUYamRPG0gx2HaILKW
wyCcPB2tgcCmtIReWpUsIJ2S3Kkc53+cdv8jYGE5d380u3pCv7K/2yhCGgVsrGGnzIk3QvI2pQgb
4h8yMsme45HlB9z3E2zMMG4mP9/LtuGwBY37GckgwZtIQiLiqDqDrNHNiP6LtljK5y8TWGg4hP39
GeZ7qUdCcT1y0/+VbjAvNlEockgV1SFgZskCD4QJcHxdD1CcDkgvB4lpTZ4AQ2a50zovvGKNCo2m
DfVEJYfrxX59FD4/sN5KbLQ8HN1Pl88qzJwRUXLbDdlFFo2Ga6LABjX5aa975rXm05SQS43Iz7Y3
lQzAK8G4mtgTsNe3TYqAIJlFPZTVMd+yuG8mxQb8+mBzRRG1eTBerAPMg3POkm6xNvaSr2LRVESu
RpP1mXMZGThfDAT4YLxBA4UhCwfSsBtmUJuRVJlx6271KMytVJxhSNwrunz47Ofql/Tk2wVpbHTf
LMPVgNeS8r2/RqqL02ApYgLCOQ2eSBKTjbIJIzHKSIciGl3VQZJzWdpJEialNYkNVUtD/eBDJb2x
8lxHb4zoLpSZ64KsdjqQqZUqDBGM5gJL9WQ5qUeMyng4sY7oeFFvKVlL9jsdRU3T5KvOs3xWQbAU
G4fPbQm2u+VCLBpm6FRMyQ4EUkWTWG4y/CN5qsB4dIRQ1UyGEsKd53qKdRgjtkT5P+a78o1Odz0k
7VlvxkZXRTZH/lyBBbQlysOnrpLu7HalmVPocZWjHLgIpbgpyH1e2nJZMGes854dcxh0Ck2E4UxC
TcyWdfAFkvCyjISER6XDpQXqwbtjF9U1MLSIBm5ZQWHzDtLnbKCR2gyW04fZC2/rDRyYaH+SiVBZ
4LKpR8aQZPKeP1rbNyrYof3dbUkf3vKaIU5duzKy7sgc7Ifo1oFhk5nKYY3WmNjjYTXgSJpYeXte
z+JZw0v6yELldxIX4rkN8MurnNzX8e5FZXKrjqeXSJRxgWSHXqNc1qBdg1xX8tzY8nyY1auX+OQt
nbh+CbgXHe2pA0HLUxkKEKJZAnOYP822siwZVViP9GlWoJNXT6PMIu+F6vZfP2SWwprOo2DLqoJV
sxnsJzeed04vjKDOIJgiLrYAwoYoRoPIDbezbOn7fVxT9LgSA+ToxchI1x8vmM4TOLCEy//87dTD
Osoci+fPg9sboDxf1OI/eNmxuP3OGSYuZab3NN23iDruGl1iHlaWpYJMQXB3zUbJrowUqQLsncEr
+q4HyMpsz6hnB0rB0cqbdatNjtVvachqHvdLolpaCKiDixRDuTsqBjcpwzP39nFIUWgzHOYuNuzY
tfv73neOn1Yl870d9c0uzetPw7NXQ3Ek0svC+SjCYwxtL9AQ/CSBPzi/Ah84iG2Evic3LTdPHDHy
X/tim6KNi0ESd4id55cttphnzQFQlIfRWD6rO3JI01lDvwBb3q6wxCq8SL6CS6HPrJmbg0YorBXd
AHB0teSGk9eCGll7gz2U/bofIaatjblazkV+PvaDZIu7UNUQuGhVldsONHCFhG8DHX0HpfTcRqPL
MDlEhQ6VkvYkVyPy7mlta9VoFO9vXDgGAf/tc58eFLnP9/lJ6ML2qK/FwnAruwNYuRb+oZ5q+DvT
pjI1g1QJk/cGGyso0fclJkiT6Fj09m/CwcxBaZ1q6WHm9fdzReNEXG0Q/yU7Z9G/ge8WljaBqHFI
JUBiZuGmqLWe7E4D/VJ5TDxfDrbV1Bb29dOD2nS51091A0DNXRnpJVgL/H+MRkUHAxpRyFsGJSBE
kK3o4dLeiXV2psEjoF5Bw5gi2dl0bm9fLAjR5Trn4KBRaSkibb9p9QyV/Av+VWaowkHK/IZlqNB5
OU8s9/3la3GIC5EKNCT8zvbvkMppFNPZRU0wEPl97E9tCBcJh2bBqfiurmIutk1bTVW7pQvoQGTU
CSb5gsABufCigT0MJTFsTG5LSsgn2+CfarOwjaAYejwzwhX/E5BAZh7IF1rXSkxnqOVriivpAd+U
vjn4cYDDMnJ2IV83L3RdVhqmj9Qmlmk/r7KHN9mNe8v2SIjITgIm/k27YrcUJE/+7sW9HdCpj+og
zKT/dgZ3cBWaHKxL9bocYoNHcIjE7mOUp5Oi5llbrqs5Wu7odoBMoDJHnC3RZWyqO80fHyN6BW/U
IWS19TzJl9UHXgL7f4fr1xssa7c0/7T8MVxgm/dstcVlJd7bT7UhSVI/6Bkj9ZmdqbT3mwa9KkcO
clWekudqhnPNcfT1Z5/CU3U040Bpfv3xTNL6GKG3Mfjryk6bOcX2tHE8sZYebIhSoHq2HZZpDCIc
TP3XTptfmo1exqtIfI5WymkbhUSzs6g8ehGqM1cJhemQ5uZCqC/ymcBkU6isYYdSBX2e92HVdmRq
K4O23TTK0vKvt1/JG7cbIxNhUqatmuVQik3NP2epwc8sZEagw8HR0DR06jCzNLqfptMqIFNt4keg
ojwA981Av4wSX78IwrJIM0fLurZaHgoZ5CBPzraX2mKv5JEPQLaLyEsu9x8vS1N4zdcnf0ClTQl+
taLql0GyoQ1X+IzItoWvL062F6LTf3RFomOPxy5VP9/gZdYw7PyHTgBph7TKgA8bPmd8Ia+Adk2E
kfxUa+q/ivxkkVXqQkFEYLjhSfKI5+qC0QwcXsMWYh/xinWX5wyWfBZbq4SwXUKrQrKfOfA1aWNc
jOxajWwoD7foj4VOo0ObkvXsLDtEZgcTc8k/GdAFkpwMNmbz1wplKLkx6RcO3f4WrW+iLoMT7Fh0
DlnGX2QZIyN2jsmbL8LCNmH2BhEhTJlw9lKLFdVfPgfCiOljzHwNFGII9ozIRTprS5JXVEpjtu9k
GQLScmgn1mDGC0qQPMiY4+AhY1kp9f4MVEAwmVMw8jM2WAhtQNTNn0eFRpCo0G5HKCd0A/Fpio9L
VzuP2LiNtX5i7uz6XVg4mTpNutHTOz+KjqzKf1+kCAEBplQuXRfGOkGwrVBR4fAE6kVKz7WigEuv
j9k+1tnOQcO7RWKjVzSlqSLhS202zmTtMCz5pFDXM4KGhs+lTaCTU4g96L2WZTKXnpMiZ2OWzvNh
Xyi+eT0tRmEwcoobFd5RVXYzRiDZGKowCKRcqIgDyy5FM+dYW57X446hlYzjITavxmdY2qr13p5z
LsVZ5eBpursQGAUdC/0DSWOfhY/xMJXt15fpsXtOhXjAxxw8b5EpnpyA0QhIrfaCU226MgU8pICg
6PRMkBd5IuMtSwjSecOQ7K4lSVL2QZ3H+EaW3jqB6uVfI7kezq5NG50rzWZ/Sh99avMMkqIekgAQ
o6S6rSCL4hKOt0SOVX2cULNkaxrC2Cyq/cHcwnbwaGylBL4Rsdc89FVFlJywf+A8f3tbCyn1lAOL
Coz40kMSSSg/rdUO/I44vvJO85JjXKbKwOgwnYRLBgROkMVryhyCkdU6Y/wFcASqwcTnZ6G/oPVY
eBJjd5J/1GQPtFAYxABEko9Hb5pH5kz5N7+aMbY4VigV4pD5ElTXge+dp7XtiBAXyKgq247gcpvs
T12FmPQ+qvK/0ykvAjGhqIUHOafY+sj4gRD7AVTHHY7h8LILY/V6ORUWQyKGT6Z5bZcqpBSLu4mc
6N+EvTYJA4TnERk1uwgaYYRhaB6IsjUXfUpVeTiSLl/AsrdhPCnEY7ymkcOeqMTnT8bUKvjmuqHV
tzIZPMu1TnCnMDPTkNtF+N40wD3ZaN/RreOMJVjiracFbanZ6GgsDb/8KSgiq9Otw3BuTYTUHr7c
GH3Mz+giuHTjjgX7ZBrtcGyZvx/wqo2oiUyk/6emP6tTLpr5fun0iRiBr6HZ/+I/tF1w0n2/PH5M
TNXsB8bZKVIsDaijuVF+7CEw8oYnaHoRgUsnS9+nI5PN+hUbQm9iE1rX1ZaCDYilBNQggyi6ZMIK
CgTc4au4/4Vfm65uPKdQvjgkGqIQXdmEOiS+4CqgCjgC6f23GsLtMMJcdISzsbSP9HWB3Z450rkK
nze+Zb2DTg1pInHVVttvt+KGNDtXwFnArOieQDluRiFZ3cuY8ATPstckAWGgqzRRV5ldBboJCGoT
Fs16wqQhkCvUDReVnMrA+5B7P5ZakvEqfA/o9s9ukhJGJUfmhXgppdt6HK7rTfDnLvHVgwBhYEae
SyUD4t70lfuhnDUszhEThViio6kGoJZ7Mhe9++dqua4mu5/BWfyJSSKNEV/G7YoTrQ8kxPgkI3ge
VwPkIWMCN1NRqpF1Oiw8n49yv/MT6r8+4j4zDOLrDiIAkLro+T9hPql5eMu2cynLNYpe0bJJO4P6
S+8jSsFBmaPElGqUqDmpGzcohKKgi+SdFW8nuvvGCtOR19fBT+RiSJrBhY/WxMiaN60AeESayd+X
v4cg0uPheTIN83tXz+R7M0GsJfl7+lLBSBn7j0HOdcw3HPpeaxb/TANMBF4OQl9ZDZVWMaqA8LK6
X6pOnKs7h60G5ZopJwWW2OQxcfKAvoz75KyTzXPLNB54XBHbRmwgrwGBEf3aFkIlnyEAJQ6TL7Fq
78fx9LZWh1/U6nJEu1smumW7FP2xefTL2b+O/Mc9TXiHWzZ7AQT7ELRtPaRjILyUTLx2mJ6x0PUK
PiDojSNbxWdhzidvpO6TzrrdLmiZwTGriGc1myYQDpWP0uMOg2YlDcR3z0wMsoUFNFfRV2hqBsaK
4YUrtQqRmhRtEpYcKQK4RJtHWBRyz21Ky+RJ12a3Heky2O7KdDo4jpJ0WfgPXjfR50AFJsFCYLaU
Zhq+gI5Hz6Lh2c3mQVBDoycesAzbOF6WepYUUFcBFjKw21onVU1mdwKosjGtNOeVYyCmDbHEiZuR
u6aHUviB0yoauvxO3yHaL9FQmnKUVHPmSGyUsJwfGrjYpNQMuiSO73Sb5+Mq8QoXKxQM5z9+xjAp
CN6BTLjAzpoWE3/sbgK58r7YAIx6ouNspetEvFZPEaj9+H/U49MxaA7+qAagdR5Rv/WkogVJ5qBd
ydUTq92c0mtUlIJulTnpXkyY1fUN1GDRjFnPqLZRUwjS7+QyIOmljfVfsuYcq2wJYKGrXVY7V487
h3Zfa8+UUcFfU3riURIvEi6xTt2HqlsyMLvMycdxYx5O0WdG+ccoZjDBg+kJ+RnLFH99E+TLByc8
xN+9s60znNtUlE/YldLTjno6cmMZYoSfRIWPvkrkt0HRkiCwTPol8xKUZAM/i2Ex2IfpFvYRrJqZ
+bPYD4bGSm0FtFdlJto7dyd9lgVsb1oUj5lOk3IHTQpvQX25ARiktY1FtTJzTcr0TFrquMJsATL0
fE3b8FqoFb3+ete/HU9dBkMtTsv4HdKqA20taM4IRu/yEcwkVp4R3foop6XsrDG1lliPPYnEb2kU
JPdQ5Zxj7P/gaScsf79y9Y+p1dzoAxOLbIXLBgDAK69g6D8MFFaX5/06bbswbnqGTebVClBWKYYE
L+7vF3IeLPL4/gHUQTS8JVlGGKbWNjVA+FGC7JHW7NQGyyhRzEDETPgaEsi6f5dg8BkhT7SnLDWR
izIYeSnbmWRYicF6QuX2Ubw8us2DK9O9+Gs3TEEJBAWMbxC797q9zNnTMAOjbD+O42d2DWOVACOD
2oups/ZgqgNyWULLLCVErS5LFFDee6w4D25qIkBzlqMnPnVCNvtN58IpEyHczQEFQD2LHQLCRB1F
Il5g6SJtp6KBor5iO7AQk7FlCpLL36p+S4albTMpG9YhzEaIHmYNh1kOhc4rOzj7U1KbmwVcJm9S
wHKsewoIJIlcPKaE9VnmAJ1GaMM737D7Qmx47otHX0xFeNEBREw0yayPIB40gay1VKtESIIxyorP
D1zGOeMfoKHp4zUvfHPyIz5Z/yPEDqSapJKY7D3C54zxJaK8kSShDnuLfb2vIML/YLldSl1XOF2T
3/irRa01hII8yEVvE2nrvJHzbfSroLtFlHJzudPeYrcYFL9Pfwc6da+9eP3yhA3lrC3X2BWDb28v
/vUxJwj2R1qOJygfJogfLjme6FzhLO46TPiFZ4aHtdXK4WjN9TUucEPYEnK6x0keYgVl6xjrgL2e
UAjPJp9TUCGS51fG+sfOF7fA6Dny0FyWCbZakcL6Mt2eQ7sIXhSTvxddn0xExbVohG+QjIWysSCX
/WwASV8U+oUrU6EPfUOOy7SINsQIBGWXfUBlScaxjnQ8H4m7TPQr1iZvQ/50gy0dn5A6sZZI514T
UQ00BycPEacih89yBCiSBKdRwJj/4blbo9SGuyImP9bl9u2doxvcM9dh9FNhouPWZKgSYO1TjIPq
62ztGsHkIZ9Rl3z9mCxYartYaTn7nVv4vNJO81+Z84/rTpLbZvu+j/AYGeAJmJSCOiU9GFlSuyZG
xqd1e0Swbj5Do+cP8IgAlo1lsQ8lF5cwnJZAjpxP6SLEuoMPv4K7D9AtmsVQeEAhHaggp6x8X+OT
Jqnxjlyb4LDmnB7JvqtexGzhJxPEiMdc64IbxhGvGIifrBjqVT5h+3VNJ4Fehy5Eg1NCudP7pAsD
0GgBxfx10p0G1ivMpOcDdsoHTmXNJDKZY6El4gOWRx1DnjBPMcEwvHdAiSE07KBd1wH9r6auNJtC
P5rwkl0WRm2PPZx9Z0cIpLlB6w+j809CafgSkBuoe9CYqYtAZvZxs23aXHat0huJ80YFvU1ApNXw
NyTHk0H2L/Wlx6v83hl6Ktys+2mxBHUenvaL+uSY1/pWDe2/34tZ8Yf8jdHhPKBpERtY3BpyfTbA
+iAh7yM1U8RW4wmIieeX9wL6coI3WDyH4CqAL2RzoRwydfSn5UTF30vVWeFvuEo8vY9MFmKcXZ7p
aVwfad67y3C3quW9j+tN4lZKE+dUQrzbP5r11BVpwBVmV3EaVcueDnqa/Wy9LUVVzTgJw5v23TOV
ex0r/Ql+bcZd1cmTfl3MwUkrZdHp8ZtAiAmqD/bBrNBByoQLYkIHs9QEYm2M78EiziTezeTmiO1R
hr7BSZ6a8pR0ydhZl0VMQxjJr6RXcCuwVuAWvc2Ws2ZTSMFNKcb4cmEwXR4xldSuNnp21fFuaG1A
NudzdTAUXP4G+aZgxFccLEeoHx7j2xe5Va0edXEfEXv3AMYdSynWLUuatVBqLrQETEWTlA+Kj1hz
mCFcPr2kIltNDIGAAfAoPHm0jRurXEAkwcoKA3ol6KZKDFpS2hkKckqwAbx2xSCwq4UT/A20w3iH
cgN49nEFSXxvCGRxKpuvPEzbui+CYpBZCnFQiiLaNYqegNeyV/vYFz5QZkQKx6gDsDMmjgn8lGYI
PBJ0X94UUeMPjVhI2T8A1OpQCI0zK+AtCfsBE0vQvGzeb9KMwBXn9nm7pwwQxQvdPpUIOWpSs9wM
WZSRYKc4pAQ1Zvs4Y+vDszWTY2PL8jrFrRnGHyW04d3yXQE51ibhk/yJ+Jy1lrDA3VUvmDDLN0by
nEbT66fb4vDuAokZdR7G6UA0hUO9lJmhqduw+zMdkg9sL/O6prdDmCdkryMRkPTIZwRDDynq0HpK
HTkH1O/HwTWRAZd0t7CztT7kcUD1XGALOndPqGdNRHFZ1u2IVSE9Ka+6l6/0d+kPaGiumww6hGaU
y1QGrNGJ2Wer6uLBgo+OetFIoDGgc4DzJMU1Bp9Pk4kequ9VvEvAeKg5x1uWzNbTRd7SJEZ0Gvjx
yWH8qB4CXWn+LHQm3003iSx+wgse2HJF0X8PeGl9kDq7Uxyg12vfy0yphGSXDdwTpV/wVgyNpOba
ogOk3CpV2ERUtXK1RGOjt5tNgdZE9J5aMP6YLmFQFvgIT6Y1+AmYPnerOw0j+1tPl9GkyJRDtbW3
8xndsKcFlg3D/Hp2ZRATmPCYHQ1+/HzjT9E4vZwX0aoreqlx2t92qpuZjFqixsN4cGGQYeBnUf9e
nkWRnt/42kwBxFI7r8Y4vRPbbW77sHetiBc045mXi3/tcrJUNXMVVYM3W7lB0zsuDrg0Asr/DeFF
lMfwO9/yHC0IlVjlkbrQK5p0Qqa2+PWiwiG5gU+OhZ1tCRlGn89PlI9ALupebqMlwv/rdjz9d9g2
ap6C31H+Nb4J9vS+vMwp/tKkc/l015kdjn0/eHWXECNOn/ZvEpYefi6CBNL7z15d7FK6rT0QWH+0
aiWSdYMLq2n/hXhxFaE5ktBEViOMx8xEyNuWE02DRQwMZY8wWPESvLpxhi20xRmj5uzdeC2qy1Jk
6OjO2iM6zzuXq0QCvM7IBFtzm0eHBRnoabY/8pL7vOAlb3Rz1RRwgwud/5xxs22SqJaYR9Mid1Hp
5XnennKQs5yOi/O+q0KkWussDu7OyXRKbtMSidZyVE/urezt8CBzPwyAWD1DZjB1Gc6/YQ87ilsP
9VNjyjhsOWLPEipmJiDq8QxPYnQCTaPtjWH6gccR3vjhIU4551TqJI0/g0K0E16FF7hVvlnUFwA4
4sGkdeS2RKXXOLW4et4iUi33zmYeB/Jg/XByEt0+tkBz3erRVqtgN14HjE09/C2xMgfhBAUzirDd
krxZ72esVItSVquUZtyFYUD0a02TNVZBzlHIwE3LVhrbcdPSNu4LWgoGZfQoHk7XahpViYyCv48o
D9MFqb1NHFoR4yx1JS0olVNhm5adQ3H/LBnn+9EKgA8mH+56j43aZoBB23ACEcyg09msmOBNi9Hk
s6TJngh0bsrSEibQ++cSxDalZpfli1t6klIKTrPle6xjI3lzhZXcVhfXJxd/Dytz18rvJpqESZco
r5ovpuWbAdZ6lhbblqrRR9GCg36AWvrgWY1/plPKtt1MfpHw6pjkhgOKbfKiyM4ixtaor9EGrs4l
WvCpLwRDyj3kBpgEHV6CW/keLgcrC9kDnaLZ3M7Vz78Lp+sJqEdVOFoMp2JJ+Ax/YZ4pgKmRNOjj
04TY+aixUy9sRYysr4UTJGYUjWZSriGuEDt+UTRLjae+eCNU0/WBx5suNL7h3M34elGnVOVoUyi/
hVX4jWj1wdrnVBXuZb2vFXGExhnj4L0tnfIBzUbo7lTYTsc3T4z9Ybji89A5TdMff9eTAeF4i/Yq
OMvCjX3W8OWacu+esYZm+0abwEjptbghsB7CYnUbjAj5d+npb1IPgPJ2xTiESsleLO+zy+7SO48O
3jhAZ64NYGbO1Cnw1HPpp+jUF9gsU3hH5B2wKENeznue/o1OoY8vJi5n69UkScjeIC3TP14OVXKR
dqQZSHjAJf3sLkvL0hErkh1QwXSXDZ2CJU2+AcJm4y42pK4ayxL1hioRqbwsGYc64r858+HZF+CN
JYMV/W4gXnEMlNm2GC4HwZbVO8KlJxHj/loJmNn3tqicASF3G+TyREtHRCLGorVILv0xraOL24hW
tSinJT8GaXEL0VHwBHMkfdd+P6kJz/3Ji5VvR23OOn7HxYoxZyDSOJ/WrGGVZh13oAiuLfT+qZf2
nNro6FPSKWflX71fVPG4qDrW27MmmwYv8uAwH69av7QL9KPzS2RFPz8KuvTwXfT4p2OZrsdAC2Fu
4jy9f9F7LfTDr3NUHLpt/MqmpeER1o1v/x+i37+Y7rwBVPpc8J+DrOhvEbr6wI4pB9HK7Fd4W+g4
c3zN1Fvcf/CVgaHytrpMB0j/0l2x1qnB6GUbRl3I729wRINmhbW+2bYN/PBX/obMmkrlEUpNqD2O
hNK88Sg7AbQ5UaDA6gAXhV1NLPK3xsnSsGF7z17AxVROyLUSUMgl1TvAoZoiTTrPeHS3isr9CdlO
1qz4wFqD+shuvsKNPEZN9+OiiWSGf2GBFmyrzFtbUfCi7GMhNaR2//tqsowBOgpWfCL3HDUdVqyZ
uzUnQweeXjGbAe9vnkxIPAeP7FgqQfTWT9NABoCI4wn6x7Eq3B63vPkw1ffsv83qbtwIR/6Qz8tV
cJ+Xg7m5xOVpVn2Mida8Uz7klgY/idL5I2mP2qtGAvuMnSncsLYguaRB69AdnUvhQBL9hIvwAf4+
ChQz7hQpoFoJFTIDcUwf3O4W8vTDC9mERk23h8yhl+1xe17GEZw1Yxh23VUQeEQnuXGsZKX/pcuq
cq5JifxPyhFMfmocis6oGfIiNEd7Zf1QpklVW+wPfR7XBB249dntdqPY0Cbfy0wJDdPZBAn1YGck
r464ndLSnc3qu8W4xtwSUqY+hzVWhP7/WqDMxJVRe74Tr93mde9Cf+B5o+y7rejBqzXIcFEfdBzI
PADQBQd+6SeDKjtfelU9YLKcZ9iKLx2nZ7yXiwYrwLTmZl9fXi+SmNcLivHSBgjMc+vieFOufFYc
WBh2m2quGaDqFkNHo6NBJ6OJWA90ipx2uZmrtEsIJZe9+awQnYAvHK3G2DmfXGv3YNPsvWiHSA00
q1S9OKKL2EMFUDx9xYtbWa1Efwv+CuZ5USeK9ZVz4ubxr23+ytS1tbEKu0irXhWV47JIAPOXhyxQ
Hy2xojieDlfvqWri/CiErpBOzfBwwVvUNbBFxMT79dGSm3dWz7v7IS8fJ6LsausICVTLOqP3zRTv
mq4hjedYfF9iP2JKGJZPHTSuMGxxRnYr3OG4M7LPzjEfAOfBlroqNRcjv3wx5vcXG6/CvLwECypk
gQA+7pPRmT8RXLZ2YtYhbi8aXxM3lgAgw2DnddwW28tS017Z8vh55A9wgmOplYrxiw8AhALAjpuD
fl7pe/MJRDCbC8iHqHAx73CZwwHaazl0ImCY15BlOj2+2efXR87eQObdCtCN+rlfccGHVGRcj0Ga
zRqx3v+3KmLzufYvrNnHCBuYwzGYXu/a2q6dqcSg8Wg9mlhd5uwxJ/54kAyDDZNCnLldjUweZE33
kq5b6fY7aO+jDHFJZQXx/pX7UiLw9kcGG+UUKBiARdnGjXXP4vLP4Hy6fLESJh3dlBA3I1P0s4HT
9gW7EdSDtte6y4n1QuhZi3HTvVfSZG3PgMEUEpJDX/KNNtnrj/jNT8IwbEqdKOOE8INpb4Z7mFlv
DJ2YH0ylrHa3n8399nEx6REVtjS2plTrMj9qCI8MZZE5hP0H0YssVo9LXnE28saMB5gbsBBY33Fn
WgHDluNh9kf3Atn3g24zSCAVBOWHJMeZv4Ph3JrfXOdkJcfAdC5e7dyOYaPyFsvlOf1qpB1HAoG7
qodGehoyhsbigwMf69oFIXvE2LLe0anYLLC2H9BGBGgToHO/3/cBheuG2f1u75XODupzLaJqfNvD
Dav6yet70A5/PbZ5PqC3ykGpRHkHGt2+ZlqnlB+qdFTKQV+ZYvrEaPtrC0k1Q+ShI5N2u0HVwTC1
LYWnD0avsKXdar4cybYz90vVXAf6dDScrWxXRJocZBF6BaKfmpqzSCtnK1Q7Qk2NcyK/c15Vr5en
PvyigO/o+io8tbzUiKa89am0DLXVzFoRMDuhckO+GA6LYOXvW+YBMtoA3F3KLsyFEu1/hhGSJSOw
ZAgrkaJYkL1JulfGh/fc6dl7AXeAMQ9kmMcjZ33H1l/MDv4XbmyQ/JssCDy2MT0Tk40TXZa9eT8B
d8NSg67fWorwDB4VZA6k9Bm8E1tLMi5DzIcnyjjEx4+COi/sObpmXWJZbrqxJgL3dgK02NxQzFSH
HbtZTVkEMlM7Tir8LJEPGtjBQ7SaHzWqNtH5fmsvZYS82W1P5p2D+83/OUTta5foaux3yCLgRaAS
5Ow0u4X/drVueDoZODueonUAxfAZJ/S9tTEzKmDJxeY3JoaRHo1RKYgMeFB/6Zi7Xsq6FhAkh6FQ
eg2LN1d2q3GR1IWtRXaB9vqlaDx0OLoD9Z7Fi5+pAJBhEDigm7ZGveAal8kKZqU56abwZPf7EcdB
ASvlv75kCCQwd/X+AFKOtQk86i5UMgwKsaAFdFH+/tt/QzPsPH3rJdE8xniraRJfWa/rxJDc8r1S
NfPIfvZaiDgrISdpZThMTqmczAhPK6dFptkDjF4HBqhH4dtp9ZqF/lFwlTnI2OUmej1DbXCGatYl
SAK/wrm0EF5nGTsJqNtwcXc4T/ZrKhnmNO2ei+BB6l6OY6O7N4oHi5usf7/wNNnLeybpRXjpl/1M
va5fMIzHQrLJMDyeCuxu1MM4awzj1Qm5f4wAtmb3BF6gn4E/ceWBdQ8ZZL0Oo4yEA5WIAYOSLPR/
+Zu9Dqugfb9BmFJDZh9n/tEehdaMFg3Ys/YP1dvPYj2FfPj+0gpbJpa5/NGRcV0m/EWH5XlSnPRg
c6U7FD4B3CTxWKtpF+eVLrdkfqdAylGUpHB7gc4lv2J+E2HOiCeALrucv0RcXmGFVCLy1bP7xGfW
vkCEH5BoyAiCXwwYhnc4ll/vypk2agEtwXOC799dYFY0A2+Hd0sASwQGVej/zth+f+cwhQ6JxQxM
nrJ/ocbQMZ653iynCH307X/Is8B0TOc+XkUyh9GWE/UEboliBqidKbgaQ4CmAp+goW1pLRzw1fC0
rnz5i8KAB6R6J9f55N7tevhWzVtyjj7nKy33zlCG6UcrVr7+rBnXIflXo/kNXw+g/SgImUkyLq9j
zyFK5J+w9QrgJZDYn3jPL5+xChrRxGXTarWNyw+Y7McUt+0KP8pryi0V1usDafpyun0d1NIVmTS2
3fvHlYkGRh4S5RpgkhYW5YM6h6725iKHNFiIT+DujyczhElqJAUmWdMf4+uWJ/C4WxOVEt9/K832
OgzmM9fHq9QJHyqpRQKSFEhLbPbbU3mOU/OABTgFqo37u92yfpYEMcaouA1St70AWqkHznZsbREk
sh9AFdRo9i7395ykpFSJEPSndXBt0C+XjO4m5xUu9jaP2lvlT+kiZxPcX+QcT4j1LwsJhyuSzbdl
QSkD72KY0TYjwl3aBlnZnizvgO7GRYLGucoj8s1bXkL4QaXREw8IwV2YOIYe5RDdWppdJ4z4LxrO
DDKGElYoNT42Qn2UhqxjhGogrQB/WsKHx6Zr6w7+btgJa/ooBsibspRPTGFRDy8fQ24rCVRfsuEO
zPp0xllQOn6FYuX+WcvRFtYBrQF2khSFeV3DaJ4cyF2DUTOJg+ez/qxLxsESYS8I7HtxCoS7/XRf
ER3Og4ADjsIcRC9OCc24IsXdegE4FZgktQqsRT1eseeHG7OLjzAaMz92WjmSkIl7UNKzX8WiDIto
1+/DC1cAqpD8U2IBUqB+zVkeepCSU3te7Xt3R/zs5oQFdj+74fUXuX/F+Adzut8C0BqvmWqTR6Ot
6atJmLfNBqp0evsuqZMn6UWgWs3ZH8Qh2EXIEj07JIqRQx1oWrq/Ot2k+VIqR6V+c1UcihAYWUbF
XGRRUqh7Kl6VC92eh/c+u9XHe5yG6vnJA/lsganXFdGEEXGAiC08fv2Rz3efDB5Af8Lvhe2uXLpR
QLmmpFjlJGIGo4fQbeMu1EF/ZxywMBifzKHzOOOknNFqmWXUpRc6cvceej4rjnKO062glM+ADxdO
d/Qu9kY6dn3+WMUfb6meFmTb3SUQQtmmQuZWufAp9VndZDMsDuLr3x4Wwl+dHGxSVvqCXL6XhgHr
fdFBMX0y85ADEd4cekOCWWEplaYggYJotIW6NPZ9WfNEk1lCB7eJ8LgCyRCS3/QxCwL3nLwSA9/C
zXdXyq/TXIy5MFb8atAmFhBG+cqEcQ+BlwefN27DgQZ51X17euhs3IPPmtzUHhoCx5QqFYJY5td8
QcbM18zD8GMmoI7qUEEDterhBYiTMrwQIj8RKTUheMskICpplyOsu57rV6ar3gE7Vzs45j35ewfM
3R+DkbuNWOa5UkrWBpr47QieF5ia6lkgPxIh23pW6mcUqeaRylLOI2eyoucek+NasXiV9hPm22Ly
LeAfsJGgG435MxdhwQ8yWY1xv0ANIvzFYmFWpK76ocvsLmHLu+7H9l3kf43DkHQloQdf5bpVA5zg
MsSp4SEN5ADMZjycLijPfKTKh6pIWjOjj8PMVJvhE+hZM9XXwKXlwgdo0eIb1vojnoTMvGIy882c
KNPSuwvRVqo9EpuXZT+dBj5UVwi5sXWF7hOgXop4goGPkUmHeFMGB+LB5Db4vp28dXLS1bdRVRST
Mzf5QLSceDx36oNo0Ter52qSwSpi78lad6Xm1MMkmSivXBxmO+fj59FZGC/r2CzDs4eLhmvk5LXn
hzJTX6kZWG8VFdCqnTqetwPStg6DgV8YaMkQ8kLoutD9xSU3I6tbnUsMsdoP7Izjk2sQq7MCG+dI
SURvN/ysZ+la0+mv30jhMW1HlndBryabxSB/TZzI4j/O++cwWpz1AJEGRqcX+jkD+es30SnZk5Vc
tXHWRAqMZ3Qcwodu0jACPn98BNOrGdvllKNe6QxIILW5/GKqrfh3dEEYs4B7WGRIDdnsxDqmAgEt
mY6316s/f9TV+kc11nrANDdyWBJCuQ2PGDNFINjTfweTWvAx0PR9P03t0xDmh9XK/rB7TrpTmcBM
CArvvaRDHRIWrCHZwJMeH5i/3+m65LqdzxxJq65jRp9EQvYOrFeTZTRrjzTdYM6aDrPajOauvk5R
aExchmHHMzHplA7H5ukmNoWIljjxfBs60gy9Eds3jlj4rKCWOXWTIXKU2u93oBVX3Xx4HEQpskLo
JsBx90Y0022jpsfAG0dp3XoI/9bZ9uHVIUK70Hdfr2bHv9GIQq3vKc3u6biUmr653ts19oVZU2qL
Cx7rVh1Eqg95AGVvN5yFqRbTR2eIa+ru50RcOXPMqW+t913qNXn0U0YtnXcqXqsm102LDPaZySlK
XZHArEG++BQPbf4oq1cmqs71hXGhrX0/sls08TVy+k7aTAcPza6eiEZI6RXpuKYWqEja4OskSHPu
iGACpTrztKJLvkSjoFpw8EpRaRwsIqX8T5UOwVzy+gv1FeZ4oRRe71FdSZUt6BGrRwHh0W/rYOT/
qy+gRJC17B7XXMxxgCHEaZfuKpsUDLtvROskrsYX9LEsaajhEz1g8bh+Ojk+pWe6bjhojkjDEn1E
6BBY5/cPm3Eh03OublfdjXoAPJcteXBw9SLjIFlwnhSJbzTblgfrxJQ7evh0AQmvwwibAmxROMXw
oJ2V5hHqH3FfAEm9hDKQnyip1OSrtDQAh1NlpIlcljA4itgAn+8Wzmt6ikDUFIlquf0LYNL432EJ
7STZMCtUnBTtcMendikObimCKYGYE+ctRqKOZOG6LjDtPssXY25R1puKBnv9mFTM4uLQ2aPbB42b
Da45f5/+MR712StXTyI3h/Xr/g/zltAi96IXrZOHuss43UHPEMgxGpeSxNd1QXl9vqrucLsCfkP6
4odsK778yJ1kWTyhRc2FGtI2moVf4lG08t07dvQwDx7bmPK6Z4D10zrSCXciQK/RPs6vzQPSQSOa
61nMil9Q6OfRIX8B2XskAmZcljMXa5FKH5vpT2GPStYL/LqQpengxVou26OoVI7LnNC0wSjIVVY8
d98HwI0Z7Tj9l9iEpq253wrFevFDjBPP2wXXV1Tx9AIEz1PA5pxQbui0w4HefYj0IOwIfzWyhs3x
6WM+AWTqDpdLX8Sq55Sbs6u15tWdRINzbEh4iljYVfW1oz3C0iq7rVUcPOheU0qsYJvzNGoqjRLv
DOr3MEx9AzaEAgniI3GVEKh1vO4O1uYqJDdNRJopy+aWu/TcnBzJyFGtAfv8foXMSI7grNTW1DlQ
DWqE8bl5DhA36M/Pe3esqh86lUjvAQ0Mn1PVGcyWUJS2YvJBbTYf85mSW7uyuJ9k33+/hrmihdjp
/N/45tmrVStgPkyE8p5VPpmnPmQSWUps4Jt51hIy/l/e0X0sAIjKcuxnVgY8LRN6yZ3gKTdpt8a5
CAtwNqbl4+DweNtR+2QgIJtKPBjtxNRcoCuyneuGOKlc5pR5Zh4l0Pr+fjYk5bpa4jQC4P9hiVZW
ApeTnTSaFeLejOgXFl3nFhPck8CGQOYI/NgcLwQ2mDg69sACy8b66rqyl9VlqkTEZCbuL28V199M
zRGa5hFZJ6G5eLmtHfX3cORzpWb5spGWJzcolRqgcZzW/E3QNJjCgFJWGzvGxTRxthTop7nYqZl5
hnFNjS/8PywrsLG6YjBBYbrXQ6dnUEOJq8BcY8pMGfngp2femebvBmRn2BcoPF+hOGtt/xTUMBQs
SvDHvFE3/GMMVUNM7+Z5mmqsQrlAuj3WqlvhlCBIJ8YJkaMwniTUQfkkXvn9v1Crf21q8sL4ec1y
mOyjcc1/lE5euUIBzwf7c+PD/ElZVTgq0HFeF4UCEGCo5ijX557qhstGBPStQRK9Jb8rzZZExggH
j3ioLFcl8rb9VmaixlmD+fW5z9hAE9Cu5+srvdxYZ76NU1leKQKKejln5RAu0FPYulojnk48pChm
AMQtCYjna3LE9RzoZutvBWOQZ4Zz3p+uFGJmD0WXVYBVs4RyQWC6gmGRqt+APwQ1Y2jV9poXgB+C
2wcCyb7KJD/HQpig4Hzvb1UH8jK/w4ki4syxQE0q2lU8SmyofnSkBfKoXtiVqzX/pN181dJ5yZxU
MMg5SWkf27p57+PSCJFIytSvAukv0H4ECmXZfZ3UUlLx2sAiEUuIuMjL7ORk+oFMZyb5LQUJJYqK
tkF7XE3Iquo+0cujpustuFh92eq2z/q7Empz0my7dQ53Qzt30wWZjWY+uM82pz2+crg3S1/8ca+w
B9XQ90g8pEFoe8D6UHeeWPc6nQbEe/28mnu61bSGELvet9mWJYLGaK/Y7ScFjy04lSKs215nL7gY
ytvOLEjvX4+XjQ8KmZLheH5kt3h6V/kYK3IaREW1EYA5FL91cLbrxoAcN7LxG1pJZ98lVKyzn/HL
JH5lNaPPHe3vrH53tEFdFZVNEWErRuz3kt4ybcIs1TPyQPZD/i8oFO1vmih3r7RWI9ISNolueSaa
/KyMtuQ1Ifpa6i9bqZPIMmnD6FljDcmJLQ/OzbIe+awJ+2sn+OlaocF2T4s8iIZj4EJFcoCuWqye
Hl7JkkW7FiqvUDLvfUzKEO0KfrNSm2bjXU2uI7xFRc9/DPqiTjv2Lplf7fy/qvKOwhqBQNMl5AUY
tAZV50ULIdSZ6athgAtlPkh6/c705o6/mYhsgtoCqdxv+/7VrxbzSyhj0ywHXsw8e9T1d53VrsbP
XJfoyO9JHuS96MqhTmHYGpkE14MuYlJYNliV3UUZUSN3T8NFv79rLxgcaTFo8IMt5J9A4zkBPXKg
ZuAnnxE6essviVnHVkHuXwVIBKfYsQ7IS7nj/xsInEKaUzj03NsuzDjSKX+DRWCmiHrf09WXjtGn
6HtW3no0mvYAtYNB5VrzFDU1fj9DZkCd5153WPao2RIaXtMWPKKlPl5lMi7uw36ddVchKFYWlK5s
unysgxSeB+Jg+SucO1FPrOYcSIVqbwxZfzb/sF6nvWRnPriS49s8NZgwde82c8HaLqyzcTg9K6uZ
J52anevIdDqPqOSH8XmF//MKdevEUeIkcH36SovIZ9oC0trIO8+KQXK7QA79E1Q3C7AK/Ozdc+hi
B/9FAHzafXD9r0tHTiY/+pv9+WmhdNqJB9GVNnTxDuJjJN1SKa/cv0EGjhf4LlhPJGse8fLt6d0w
mqEd6zGYwEON7ZDV3KKKVBtuMqcXAmbLG3cepfn93lDhaqB7ZcfytbRHtan4UAXRQFzVZNyjp25/
bBVTW8FT87wWisywxmrPU7zAoQuT/a5jOShnf5rdeYawc5VSsarYAgDisrE4VemcTKFTbPCdawZf
LxdKCY5F+m7gQF1wnfd2UtGCpqUbuhBFxv3xO+9P8T+ihjqX61S35/Noi3DVGEF7gSWWVfm5qlUv
kK7QLnik17ST+/TJhwn0yXp17lQXbvT3gHiP9EpnNfFf299ZH84wX+XSQ99XTqAV/1JC7zUAEtae
U09CGW3rjDhfNTHBWcGjMeT6yXFrZ5uqMcgbZxDA/g4yxdtyzhA9PyBwsyFiXecJh6DrwNUWwo5W
kXklTVnDJK0rWC6R57xltjqHVc16MfL5yBgvr+smIIhRcm0SAtkrerCBO/U4RFlCe5SntIOg7cnI
HYNRoxvEY3kBL1SQMLCtPpmd1SWA8Fr5G51AsbekCVcgjAAhTWcDK7qqlwx3vFxKCRT6ZBxPQ5eD
iYyI72u6AIayGENLFFZSU8JLus82MSycpAkufGmOIfvGOfP8HtCAtOqHRxl0rOHa6yJGxo7Vc7Pj
5vWhH+gi9339qBWloshZYYW4Bbdofk9sHGF88sXQpzUJpmoOKmFylFXMW3CwnEDKPmU3qcCR6h2s
sExKC6CCVqKCa2B0L7FK51tL56rKPxLHR13XMo/SR9JSzdCH9Z+ErGM/pPafRN/o3sXd/sPMVERt
QxwJiTs9kzcex2a6PyjXZgf4d1E8A3udt1vXfFgtUH6e4EOJNIP7Iug/5hfg+sQqmEvk6NDFYwq1
JxYG3oWEiHZp4OFjaQPMY3xc9s+epYSb21LN1jX8N98fte4okexWN8OmRJIQvDrDQQy/7s70o3xH
TlIeuF3ETJTIpHlWxuzbuZGiN5FTZNvrvpzb8Ev/hKyTCs518zbuoNUzmAuraKkWtbqebv2w/lnU
W562LgwYh89VYStX0+/JwMtr60kbOxz1000gZsBo0FHaXYeyq6+gI2pddbQh3fBXmV6kcZelgw0W
hdrlS+zZAkV08YSJTKaYNt5lNGXnnbCjvpVsl+c4jlLwTp6uwtZaSJ6gtU6mISrVqNd/DyXyTuxN
awk9g40CRJyZs/n8SIMUOjVHodlp65a/uArvwyeNbuhzO1wGsXmn5KVFdUKQE63U8RfPSvZxTeJl
+pz6R4NDNSut8iDrmKUtz4Wuwt0Zq4bTJ4Z8v7GyUTqFoIXNk99uZZH9kVzthxMDFP7SgzxuTcV4
MmYXTwmbGnCrbTixRBx+e95Qw95Izbkrgi5/5fL5cZqvR51WfXiRHVT45rlgWtbkySc5ZRDmD8jU
Ptsm+xiMwlIdRfB0YnBKIJTeGgG25EQZBjbzczFUvrUBQJEklrlSsIjA1nZRfXrr6e0DJQYIP188
0G1RDKKVkG3Z8DgSu/nGP7T6Z8qAbJl9cGmFwY13cO49V2jkmAybDdR3XESFO/TmiExeClRBXlEV
recibRRHlclkaex6otjOePRnbj8HW253giOFDI3YoqofdBzZVl6ppe9ZLPrCJ7RJT7yaMODZeJn5
v3GPbqvzC5HItnEMksx5eNjBpDI0LVCtzY1vtnVCGHswhYt4/x0ruAKVd42cyjrkFZg4/gXG0Dpe
vKJid20MoBGiP7UQ8MK0vOcUr7mdNN/p2b2/LvoVPfw7Ks7+tIxdgVRNSkaNjA+8ci9Ag+JiweBI
m3prrtpiVFe4Ci8YA+WCO6en1e6aFR9KNVYLA5lsit3BE4+P7FWtWvs+QadLoxK7CJfNTz4eBoBY
WM8qgIejh+7UXNkm+gMNBT3JMZhEy7hxw3azqRASzytaDyqB9Fj/MXeWr5U97WbIQCEb76V4oHHb
P0e/6qQpFN+f8P4KnbHKXCoxRkJJy8JwyQT8smAfbT7xS2DpjYHgA64tnWT7BCjV8MXXXr1HVJMO
LQwJP+tm+qH7OliL2BbOKW1F+6rhrFCi+eMnEWjIS6Xzb2cEcWeLEj761JT7LFn+w5pF6KJkMlny
QQDMNT8+9Hp9Ue4mWbc50iycuCb85Gs5b8aj/DnQNbV4HCAi0Zk3F7eNwEpAXRIs4qY9ydAEUoau
FHbzgDm4fYJjLibZHyZgC/lTBX3GeHSc7P63quU8BphH+UulQHvrs+KO89GTj60mLxUq+UP+JSiV
jUPGQwLCEs0DIr4ExCXcFxnT0bFYNYrA33M3qPG2PEfhgEzO7FBRPeEtM4t6OEejeJJgHMjFtMdf
/wWD3AVCwSGJ49et1npXivrHiNy6wIJbQ3W4GEmOPaUOK92rYvHd83Zb2sIGrPXxBPRhREMWRFmM
Qd3PAcPiq0TuFhvYUlYSCtgniy+GOspc2F0ii/w+6BL8YZlUYzGXGjdV1kLUIO/81GcsvvzbeAoF
dZAPewJV8Tyw+pcT+8RsBlK7qMdRXmnopsYqlnjh7b3P2xjrZGn59uFnAUyaMo7nB0sbyjwg2qxG
PefFvmnUSN+ZJ6F0q4+d0kwQNtKjawehQh5g03gzVBDDD+Vr7vSfPfORnNcxtLyWTusKw6L06Vjk
cTt8EOFirDP9X7fRMcDSl7KQIrI9TLLMKFjmMj1Z9ojG1RleeuzWOJ4XYFZZoiO/N/X6YUGgdTZf
HC57dxv4zVhC5o4AuscYkvVPOu7gD6Dr3smFPJmPMoLePQK/Y2S6ZLfOPKmANbM7nNhsqios959b
Fh2J40V2SGrfmtKYb8BHG2VpmJFgiLi/cIF8sk74KqgnCEkFfaCLNX4LkiEAFr2tBt98XR1UDHzY
VrzEYXbkxjdZLcPCDhD9u6cacoePDZK55cC/wtcRIoysmh87OGIui6XJhe0XwEije3G/oQLs1h5b
OwO029tczLaXYx/g5NXqGu2pdgzoWml8+ISZ85NvRbVTm6kpu98WsOzZ0E5Ns4lZQASqW0SwHiHI
oTqzP2HUzcctPxRsJ/EnaXHNFqieBCHgisoT3wXrp+6wceFti+N3iGGZjnwr7g185m3xntOyv1cb
GfQOqTAze1cuIr0iGocmiYcVU1nYQ2e8y0JpFUWp/tKWJGDYxjyJuJjho+g94fD1Mcml5qQEUxnD
kNzKik2R6HepINppZzf34p5pMUhZLPMHC22Z+OJVyQ9wB5/roqtrNoj+sDbHpJVVktfd5PflWUWe
vWW3PYacTCxR+TQgDhPrsxk0n8oMNH8vNvqP/DtzlbKOFrJlW3kihGEiT8bMYYw1V+EGdE/Up9JC
eUe66YQiQk2JLJQRNO8kP8Jvryi9PV/eG0nkmZKT8iCen+8WC08hWp3hAPftQpR8fgUyUKIKCztq
Q5jvNVxNZl+unY5ECcvX14oWwA/jgbnFjYn3TKg63GiOp9CkeVaOpjbjn3F7GArDI3gnQJRRmrVd
aPyeOj4phaIlg8kU9nyHIxDA1ns5ZMCjlGjwZa5SxLHGTPysmeDQ8c+bmsL6X5+qJVH5pOuiViio
Qh7nHtZd5gREYlXNOPpPy0UGdWhxBLfrxvygCxfnKXCaKFhc7E/o73L2FfptnUOpV32d2c7mmYp1
4VYNSK2cTlYgxKBz/amTO4xCF9sRQQUQWA4SvosTQOmiOdTVi2pO0N6lGKQnVAl6mgKmVfIoGlJd
GMIXPI7exoL+nSCpc0toeC91IOAYZqK4Zn27isVZ6C4V3zyszIz0cUlNaY0JsvH6L3wFAp5W4Zn6
nNBvCIJxDzTusWLqHTdCrLfPQYpjFjpYlJOq2RFvEq2B3f0NUS+RpPg4qbWcSD/xAoYX9pqzjuMY
yuVGFNRNTf3djD9twggyBuHyss06Xm1KxkaMn8SKGGOeeJW+gsZAeWf4Db7fCPUWgpL4Gcsjhi/b
Zbj+zRHifAoRqr9E236KaGzJ4hRZ6S56d3Li03W18Apif/OM6kxUskddoe/n9h1MHLGuT/ECmDvB
ISe8wRMxWB4EKvdu+4GPkfP1ADLaUpLW24c3slDfpWo91KtYoUG3CDzXgrKpi0XcQTZ8IfxzJT4n
o6SyYEjad/D0smL2r6tUq6Lo1/Eti/RXesvE2EWMkrQcI7l7pdK+e7+UXVMabADgeaKIk9dRaXr3
une4BCBfxz/uUTb+e0HD5L1Rpv0JLmvE1vlFeZYSUCctvwd6tGbxd2n6HNCSB+R6cK7Q1nyckamf
AMAqNp5c66gUXTTtfwuXSxb6AbHW3mMiK19Lbj8lQzia9v7ycXekQ1NVJW4LCHl36ApVtKROO6/x
Lxds5cZ0IIT8W2xESZPLaL54m+8HAQ3cWxQ88X8wgIHZxtsCPGgUEPWP5O5LFK0EirZgRZ44lozd
nAg1nclxRf6uMoeKKctQeIjycIfMrFIMg2d3CTrKAJvaK14UD+AzIsjFjUhuaGenOPL5B6jyGHIE
xtPUX0ET63xkrOwO3s40Y9Kil+CSxvU5YXn19raclkjqBpJrezW2QkPkrLcpHlRn9D9cqT4qY+p2
IkMq1KlS5/F/KRKo0QhuskAn86XhDHEr+1feSMF8SxTGzo4YGaaA/ZQvvgTohZ5V+CQOESjtWHRB
CmFUGD7zH69OfCJafuBvtHTFgl6CCt909Lkz2KMb1Vou/2p5pE+gP4Y8tH3l0TF/MYQGNDW2wPSM
7wTuAIPipvusumq2UEbBxnymGPo75g6QUYH8fJ2IK5cO2cbWgDFN6DVXAUXOpUn42TEOS+GV9Pdf
NfjW4Nr8h4S6GnKfm9aBWfg1VPVfodDvkyMNZxNog+nVM+rBp0VqPzx2mi1mZI6NU3J1LPN5KcEj
TLvtLgvH7I7wbn89fK1Zsp6uUlpbh4f6JzhzZpNK9JB52kl29ciUuHk83bW7r8f97dXhfAZ9Scf1
9G+hWQ/fdK4osF5NfF2EYeSUCwFSst7ID5acj1RhVNsVBuB1pGNYPNbftIN7zwBWgQlpYNEO3lSj
e68mXWWs2hQWtmvoXnGK/3h5DdoxFCHcwQdDTiU/n+dc0TXQ5vVHTXDAgaKG0wi6QFP8WCkSysRF
smEJWftOXgLtAIpndLYY+bw10TtxxReoNo6GDaF9/2LP3jov1uEMH6zEtjVOZqvd4wi9ko2y8XVU
y0OLeQtxsgaOmKndVFv5+1V2ljE2YrtR0wZSclTKVT69mAIkbhzOT/nWifMgjcBoG+hmHEFgNUsM
3XkQUgWoq2fbWIWglGmKS2625VetyKNXEzYyKoc+WzGhQuZJ8/0xSEuOVSSIe6AYPP8K7k5/KJc2
xDpRt8GDVsiwesMSse5RfKljjfur6AuRidZJrCFXNlPoR0cs9+TkjltB1ZxWellmRtsO4PZsC2qg
PvCzCiBarKWjLGLS5S0ONYm+wDlEsMFzLg6wWVCbqQrfLIUL/J7+HYscMrVmBmK2GJs13IGOkTlz
gkxTbIhsV/S4hV9t3XBHM/87ReTFjpu9q1Ta3bZbjMSqTAmnprqxXbcbfs0MYj18xdeMQkWsUSNX
Zh+ivSPw/pLCVHzQCGzARap6dSSyOL4aIAFptfOlndCN2XBWhNn8/BAEExFrtQVB5hmoHXvmwp4j
OWXSK77NXqSHF4WuuOGjLpfbv0kVtXMp80+xpo0Xh1ukpKmtckJ5xzyItIvXGI56l8Vyios4VUyv
H0monktpzqZUQ7hCxIGkIBQCH+P428jw2aqYnEs4g03LH7nMYHmSirXQGdeClWTwt0Y4gRI5oR3Y
I92w4l8VgsaGGxlu2PrEePGkgalA9REvcWuPSf91iU3Pl+FG7JH2SalmP3d9KD3nLzdudKkoHwmx
FEbtTqC2aX4abrWAxdZv2cQUcB8cIn/OFFpxKXJjv+tDVcuH7iaLwcJ7ByX7y6vDsscaZCrHKGxk
lSJSJ8yBp/6sfMrwNqquZPOPA4x6ltIxMdCdUKmVoO7GnPOtWKaHqH3xSLDHwzzk15zwknPU/OMD
z2A8YE6J4SFBNWhzMy6rJ4lIQfL8u2drXnulDlmkCwKEebZ8ybDbmth8aZIxyPHKSI6PVUVD4TFm
DwsoQzBRRsOPy+h+EWqwEMw51HTGYJGeS9uabMnNdjA043RAtENhk98sOYCpBUu5Bipe53OEsFMQ
CSPWg2l449uNxphvEsboAiSKupiju+vQNtUhEJ18Cdpr3hS8gz4q6Z39YUO88M6gtJxdmB0LyJIZ
MmPXn1IeVHKrS6nEEXlnGhhFq0LWWpr2/cvZSjf33FpmFwKnehLAnI9pgwMjWPZ0rBriLn6CC7Uj
JmbRH09iQZXuqkN0eWlHXh8aI3mfnPcvHEEvpCBGVahSS1pHrNWg5y3H8/DFfE9AnqeqWMi3Z0pY
2v94gLtf3opcsy3ffs+bG55BxJeEGbPEZj4KKt13InaFCGcYfrH1wq3x+Dq2bHtEcX7QKs6sT4PK
67o0ZpNHXBkmgM8V4L5o4GxVKf3zOU4dFn3qbmfDCtlQuAVwT1HtZY+lrOJMnHOOmmfAFgV20Zpa
HbHIIl6FkNMY85RClSVa40xMBuWZKMw3wmCyiBEo8LZtVrl47I0b/jBUC9f4vxo87tM9oSQPN2zV
9fqOOTHrvInTMMCCIxISD4AGlpvxEzGm2Aby+8z5FrYdLW8VN08DNN1EtVyBGsxirILVNFLWY7Ez
7/F7fdWnx2fUhvmyWWdy+Itp8Eq5VJEaiys9s5q2OX7N9RTjaXQpQDGM6ED9NlWxRomP/gQA4Ddb
AEj9FXkRZEbLtFpqyNBBFpaAVUttjxtnGjMlQ/LNXGscSXVd94VOeJbAwXDsd295pX4C5rf/boXV
pzqRc98hP2y8I5iyI0ryjC3CBjmesEWEaw9nkssGK+lTGCQr8TE/x4NRVvhigcWqIwNp7nCeS+zO
lkJW2w5h3tGDnKyocfJ10t3Ij/EgH+sK8B2gstRH1M5kNWpyEZvwfLBznyjH/Mq7xT66ztV7gqaT
fCintsfuAIpngFVsUp/wEnYr72IwQNoqIKqlA7jY/CsFTVT9pIdD2770rFvDwapY7bIunmFmfysn
yfeY70EbZCP5y1dyXVHGnQNHV0Vv+cWIS5vQJN3xho3HE5L5qoj/+cxT/gGkPpeBTd2wscJ992w2
eXzkAmfxc6jaJk9wMCpL7yDjCs5ge0urYYkNy3dUtKuCWJxxLXMeNq26I1sM8h4Ty3Kb3w5YqC72
0uOALx7p3quK7p9C9D0BTVgXfyvbiLyytPL0w1ldFKLnmiPJNZJCtU9e0QoqD4I29sdCNndb85ML
PTKkci4J56JBAmWDvmRC+FkqP83+r/zhBqUjLodYwgEG1fBLqacMjN5or0DLEI/0vXCy5ep86M6i
UR4uQL/wXjAOg9UuDvEMAO+YF98WYPKEng1//g6VfVriKlHzKVp8uzEn6CUWLi8a/w+5vutAfw2u
3TfAvFkY7Y5mp1a7MUmJUfE2u6MJr8R03L+IIcqtKXhj3dGaUhXgfVo2GjoWsuoKiYeKo04q3KwH
BY7XPhoIeuQ/ZHNRutmJABkmF5L22Qd5AERB/yzinOzquUdUUIsv8+KZGYp9gsKmGf5JcaOAIVcs
+Hls6g5vFtRlweWzqlNqknQrOjKmgcnjxrqnRa/xbUKW6daPwa+r2Ujn9fBXjkgpxctmMEbd3fXT
34hGL8GjMi5h88ACmdHPLUU0hAWT4LozrxjH0+qPZu+z5E2luq5F2RTUehNEdzilt5bC5QEGrOXd
01K4HKQ24eBZnyr8+sgMvodotydDcPSnjdpzcOhzJUej1PY8QnersS+rH4aD/2LoAWf2ZmdekvcW
F+mi4Zik2SZdJCUDG/7p2zF1Pg3JhQAFHzoBEWtf2XDC/ID1PriAoBBEf1thkvrUdsgHVBImVxmS
3VThIOAVFeTGK74hCojpWzxw9fpk8gCV4Rkm4YuSfYytKQxWxO4KWTumwdLg6/+JbhOPLm9OPf+f
hK9WLM6M9cPNPC0+bLXeYQ32pbk27X0HZZKOvMm7UlhAHNuKMhg15BCx1yrL8ySffFBm2WK24TjM
a/aq6PQgzNWk44APvQ8KPQ28Lj8LGGnuC/GagDcVr+U2xZrE/QDguNU53DOsjzrE7d5upy4XrP9l
t7dlzvxXT8oauOjc1uA5aS7niHWsoP8eeUYd1GFTOurO90zyrwUayrzIrtjo+bvXndRhMNAZmOij
dZT+kgou8JQAD1IARtwqpYJD4D34rZSZHyqxLW017Teyf9tlDBNvuZyCuAOddOgCoVU0G7BcqAfA
iCgw0BKy0mIBDSM6t+HMvtUwOy5XuMPWXxkx5tky8Bh4XIEBPh6cXbHHFURs1fkJpacqHiVBdMbl
V4qjkdR27Y11ZsyTGY8+2epdarBtYSP/qrsDQrZ8XOrRK28tM5LGEiYTEK/9zh5OIyugFQvfEZZu
ZXmb/RsLUjVvhhlnysNCcI1LuEOjLr4xTV2xeZQcw0l3LICURil15IpDhXgv25D1h9ivlyhfLUgR
0HhItT+FTdDVWRQpt7iqnmlxzoNdwinCXMj4GFOpC1687PwHDp/VbjTsyeCU9uAkQgrlV2vKaeTh
uvo3uU8ssDypM00KgkNePDpIZ+G3FK3ngMnhcg7h5UiJXp3higp4wnyxRgaGcRisNdBOTYUn6W58
FDcVphxbPRs+vA/nh2PnwJ0RovYnIxFFMWEN1hxCouj+Hk0yEghJvxGSP0q7XXXY9x373AExhd7f
C9q7W4Wr+eGer39cgzwXhrWaPlQQWYvCEy8kxbt23f4UPw4bhnICd5BqQu3oSQlgJTg4EGE7/31a
zdH59yluJmaTTjGg5ssks3C6N2sw9WjZZDZI/bAaz/2bV/RyeSb3BYtVxHw03F+d2hq444dkM5ML
wmYxbcfJPY3kJubodS5rFQs4z2KMZFbpTI+C67N087ZfH64hokm8x6WF/WdnTitWpwtCHhZ8O/VL
Y0xNU1ry4o40JOIpsc5HFRzeg5OupzFQmiwH3k9PK7gGVpKcb8S0cHaRiEjy/pvtGQd6rj+ollKj
rCkAHT1RQDxeXPcSIfyoKR46lO1O0lK+aNYzCpp69BGk5CXezG6hJUoiLbEbTvVMMXFDqOv+RmBm
tf3FnDDLEvQDGeLPNGEAL2t6R6JqXV8bPMItvknmDq94ArGRgNesbQ0Aa5NewngvG8oVzgMI+wqS
5680VzN8IYD2Y3GZgw8/jel2k46IfUYL2xE37J7sIZr2a0SVcJStaAiHzTVuf7DoT9UR109HfYaF
j1ERtu0kBfsTCX0Rs8183dVF1ZhXdKMtV/sXiyIEivsylQ88OXBxKGyFBFbe4slKqdp9AX0JaI6W
Aykxkz8QBAna/Oys9FXjzylds217y99pWbHPprGTD0wBIFGjpWSajsjU7HIAHFEk3QF8Lw10sZ4E
l9dSISCcQVs6DTVTTdXfIVuR0ee6+LvxxMi2Q7kGHaCLQhn2UKtx1qIzBKZBYbFVCdjMBm/Vvv/O
Lrp+CtuMYeL2faTUVJ0BnODNP4R7tQAbSAat77p1Euw9HlYTiboOs6PjRkHOidlzyfCpvAZXb9Nm
FvafKz48q9ut+zfadxOP7MH6Cf/bsHGD+EYHCRLK2SMYTkcbqluKTGEy+eF0yt8U4wvz0lQeNKvA
z0FzYZm8RALJfO+7bS66bDQOXZPWRnzfVtr3n5CCc4vtCs9xjmVfbbSnVUjzp4UpbxMDD5tGxCe7
J2LpJn41GdsLXN24breuciiME45rwN9txSvTauWFkUHRrsk20euTvdIag+Mgb0cKMmAsJwKmQpxR
Y4y54uEmXpDjMWH3LkRZKwNWPrv+QoXIqnkcv19ebR0iF92YXTAysziolX/NDbX26FU9njNLsUn1
t/Ho7sdnCoYkB1T7Eu6CfGVjjgx3mlwkLqIlrv/Hyc4f7RCf8ieW7hph1gbS5mhYgtYe7b+E0dQp
ibrLCcjDPV5W6o9rBwZ8nFnmCL1UWoHD409lM3kQ4lLkEYSK0coEvnZYo384pF+ZzQUI8o0SH75O
5zFaiuk5ip5VcLHNJxOwIb72Gyz/kJOuK7k9fd1Hse5GPIvaI1mU05QW8xM0GMGMZQsMn5AKhAmX
AcL8s/8xgpOkLStkXwpdD+R+U3HIWl8CLw4t/vjxOsB+euiqJ8lvVbTjkk+KXcH39BhOO1IPqBiD
Yabn6kXDJ3CaZqi47IWJcthu/KnMA4l10FVEdRkuhFuevsYLzC6wO3Yguc3/55PIkBZdoxM2hsHI
OJN6eMm1u964f0d/xBq+kC8IejqEXsyFv6Zl3do4FLW7P9AofDy3NVsZut5YKItVePL+S7kLBS+u
4HXoYavFAoREF8IcDFF0UhwUfAnDiv6dRIkDAWlgss6hNDMQ+eVgidkKRvxfkwbncueGMnXdZyzg
EcDB/TscNHwCIGxbCuHibXwrjBP31AKIk8apv85ELgAEzkrRcnxTVweetmVIPoFwSzM3LBbONpmB
uYk9Ln4ivKwvkxF6t+VSue5WjUGlZVkreU4196DfNsmDLwIDTNerBj+ok6hTnuC7/9riV/XW74PI
wLIjW9+Hzhh7wOr4vgcoWva6KxKMl0+MxNc9itXt0xnpdnaj8Oxac/77D0/bJbgueZ6TAD0IBbmg
JVGtXNefkZeS2u1CnBPiwXPW060v3/UtCjdVB7dJLbVuJs7Eidnf7hDpTHncdfSYrkFfIcVJ6GcP
NNNoyWEeqAlTUuHxb0wUvMFZFeKLmbG6qz/5LFcFagY6euHmXcu3Y5zC3dXzlwIy1MlYbHZjvB35
95srXuubnhdDdzmFQ+9EXEt14GrvIhat+bJpaOAO3M9n2WgscGvdGzDD1EgsBl3d4vj91XBga8KU
ytRF4VKo35/2chrgMEoWCVEEH+ZsR4alDsmoJk4zSsbH0QqGDipnlyUtHsgKwMLaeR+PlCrx6RTZ
wP7XSCAg7r3T2GHpqdlendRybJPi7/f429fycG1nJqTwkwxk/nyvBh9DOTP3MoZ5lwkTs6MsWsKK
PlqvxPuUFUY4KmQDNSp6ceDalsxcJnNli6A77FyAnQNQNis/QXHGCpIGSJ2kJP5fI1V2vy3EKxma
1aC7K4UEeRFeLPRSIzEhYmJFJTnI0d8FMCLJH/hUZSqr8vVcAOJQ57A/CcmnqAwRZBStKFFmujah
WLCGb3vuQKD/pYzalpNseekgWvN5+z/gfaRnk4yHuzKT4W3+4GYQud8i9Y6SOFFx+9iEOPQk/IrL
SBaPRVQXX4wfnIE/CagztqhRjgosmsnM0SIHIMJMZ3ej1O9XFJBB2nVVrxCHImn4me+3Sjp3jXQH
kpAwE5m+l0UPYNkX7HboStPP79i/JiTvWw3jVR0Wqn4gtOoNJFtn8CHZcVKS3zhcAFODA6GianSl
8gzN4/MTbtN71xRBadZkMLpgDbK+XwVmqyYPP5chFITNqHUEj02bTB1/RCnFGXj3sGKqJ/q7tGd/
9CyPA1XB9iyHvlwZEovY2iJ/yBk++YhUreS6jxN3/Yi4SPyEhpWDTFi34q/PLxioMAmhAdRMsVFc
/rLgM/NuWhwAmJwCI29T4abbm2q2BHgZifLTZEiciL3LuDR00OoYTmsZwIzu6bbe7p4BjbEL/jYK
qmtwDf7208Izj1dv21Hx2keg4b49v8GzjKTl5btPstSqhJcM4OBm6IIe2rYrknb/n3aqPHYckfI3
EFXVom3gbrYDD1hdyGBlahPRXCJoIaLxhx3MH8VJZrZkFDE0Yipb78fywq12t+y04n2gM9jUmOyb
YIiXSSPyPYqp8QbAxonycefY7i+TmyQdxg4JqyYh+lRpxGW+c3jHgGEtD5YYQRCNmI/R+n6ywca6
pcHFINAfCejb/F3dqjs0+JSs+LQOtAlyYRPluhRwOCXMNYnwqbNxBkXQ96Jw23oO6m9+ivXwES1b
tHczgV5pWfiqxzK18TjL617NvIdyu+vqVI4nSENtEr/kecQdkJ3Yw8knLT8mj7B8kPa50xb9XV02
VPru4M3Dvo2DvdKN468Nu27fcd1fe4NBTfPmxIgRs8Mezfl/UYPy+hQWfhTK+/TQnB6GKE45F9CJ
OjXWlZjQds8F7Wiw6hTPs4YGcu026vu/3yOB240L9tDm91GMEUeiM2MdVwbHSbDnWrUcXt1LJdBr
+pckzL0o8vvQ+SUkGBcSq8sMh1lDIbizT8LjgiLlk/J/PGNsUm2tgAVchqct/zkbCoM8v1/3ImQK
WQuAFXPRc5k2/1QujA2OvHJ3p0oiWEYW7mS5sTgfbOxr+YjJhZb476OGJGYQK8gH87i5e6ZZTEKE
AVunHZC3AZpZQZ85IvzQpEDQ0hbPfc+wfBogL+9gzM244ptumsd7Mm9U076/wZZx/cVj+xFhl9EZ
3iqBdNLeLNMMv9ji/ndlMR5qjbHeo/CqunqEY20urjpTaPgDzGEyMLFxVRLcFFUD1eGdDUWKLfEr
d8JlU9043Nj4u3KLveCUx++EKHqxrVhYeE4tMWBTJudQ4DnGQHMy5ILeg7AWIq77OGnzlwDiBc6p
GgXnbNcV3Wy+GrImLhIT4O2e9MbI2zfw0JLpQoxQLP8GOi5XzwPvriyZM2utMZfxwcEX97AQbM9q
y4Ia0C2OeDY9YvmyDSyBYt2Foxvfkhy/6+qQbtsNH8/q2iVg56A0Q6lnZnWEhR92yGQvjpd20zFm
OxWRbdfMoOJwRPNHj3EXyOevjwpycOUwosSgBgKPloQXVKKpXgozL5cJUdE+P/db5Zb7m5rqhdm/
4/e6BEkmLcbRBO1xJYUVW8tWZfqsbSuc6deDp/EK42sNQZCyNbCwhMmSoB1kdgeVulwa9SMAOw0H
uAudIBbQOHTaT/abjMzFcKn8fzWEYePqRHqlaynJv4Hmmp4a1IaIJrKTnPJ1ZNN93i7UG1CA4FxP
ATYfLZtuWLxNRkc1q+aFz9p98sM8jWi9utqqO997oA57Mx8EEkEoLhbzgLdFQGrP/uayIouTcTC9
Enlw5VIFcAWkS2vFnrIu0EEg/RsNgOc+5W6H9CAsiHPRGcyA8I9Ph/+YKGinf5IPpMSNTRB/X8rv
d0t5qnOhNQ2MT0CD1eSfGKuHsrGnxnwgVIwOg+rH2CzgyyY/JjNCsD7ed1DT+GuAYi/ftWcaknlA
dJeLGNqMf7zcf5BA+to5pYgjU7B/YRDOTx0zPfGTdVUMbEhHu9eatAOe+r0NdHRJqUCNg9mHDr5d
PB8rg7p3+TxFOdqwAJSaCsLMY9ahWO5kJVCvVQN2iVA6t+1qusqnEjYTAHqw80BnqrGRGp/9QnHq
IzgGcD2oB4hd72cHH7Cysl5P8mB1E1EcMmHS185fWRf9FCNcEebz7ZBiYwyfm6nmzyArZFjdMiSM
0ea/rlkgr5yrwPNaRroTaKclC0xL7BBllTx9a/Roc794OCYHW9074qhZgDbG5PI+5zrOSsgJTenq
50Vsvnj/XoNC3s2uFuMrbkN7z2N7q3Q2yxibVztADU6kzPLoMrWDCF5u6aZWFe5izGmj10qWSGkL
6jZfjOt/0uzgrQ5TwPzkyE7ReKHoG/wk4gOLPdzM/ON+YCVMMmGIx6sZdFGE79disxydl4vl8apF
kzGxU7JJSyFhZ0N9TupqA/ZX8ab3+kNx+EnCYfPiFbhFcAlUyVewgz4H9y2xMUgucxwGZGgSupEC
y6lEo9IyT9yKZg0+kTYRAp5tv4Mzsvpd8WhkdyM/YPgQe9IUhtT7EBFxa+IegTfZQeYc6PVx4K1Y
xL6G1JUp8Hs6agtZuH1B3CPeNIptT6OQFurOgWEsYDE1oL/QGaWMWRmDySqMhYMAAzIj49kdQh1p
caSOOlf51QsRPwjhejuntGJYb+TUpZ8SW1etALNo4XSXeE9hPxZThlAg9TTgDCPP2w5xYRcu6L4N
pmnxMALU6svpdKFrSLWcWOsmzHlGrh6dL1ptl/v+fXzQQBxEXwRR11WZynUaMCz27vbahICkWC1y
n2wuHF8NfZLfqBcGDLos/nyL+p3+88kK35xvJBVf6PKvREOdik1vH60OPe88QN5vkScUkXpSEqQR
JDUKW7BtZfSM8J4Ufz1OIIx3uLbE0OH/2pUC8xgRUU1TdOVN4NlMyapwZK/Nuw2qJ9axnFrX524S
hN2acNQqJY9MdhGDOWr1Fr0A8+OAUFdrunr0hj51PVbgk9PWCiKd/5xxhCaunIIYNPV2lVwVRO24
f+PCsX377wVvCBuBeh2SzORceRpiyypvpJHhEdxjiRI3hK1uAWc1ee5KKzE8H4YvpMPeHJH/W41i
2vxFjI4F33koEKOpmp1xQylxszDd8yFQdJ0dq5pXg+/UFrwvYuhOr/Xt9se9tvF1ZXxZ3/9cfp6B
jyDtJ3AzxlB+Bso6BR23jp/+RXynn82sbjJn6LP/J9AYoBXtezV0HYCLedXLJTZII+zZ2XC68BLe
UlrE0OHDsWR1tRn3MmrsvinhD3VAI0pjheBW0F7N5RT3wvi+UwA+i5qfN+8UzNF8UE99gp9R5q04
apiwFFY2pDEEUgRYg+Xhl1aYVz0uPbGAk6NmpDrgr9sENjrIO83QqNYZSjYT5ktCC6hHYso19zht
Y4czeKGucUJwsA0XQoCBj0xNxYdOFIse7BVrpo8C5l8hqCuuVH5yJt8ISXB2xPSLquRilRbhfEvX
WyuJHLl2TOTptwQoyHvguP0tpRU6pwdDZGFgFvx/7IsQ0+6rcOWGDI8v4639lpW0OrXte7KmAPTG
PXZZ9lP3vlYCzisoB/FTPFTQFlCQnl15p0onEyexkEbYtHs8Y542lXAPFdJGASfa5rt7zSzSWZsj
V+NqOYWpJXBwhSzk5kS38skk4/VIwdkuFXBPugOLxeo0/vfy7ml8PNvS8RwEcoP57h5v36SHsifN
YrLmC4wzA3rPheH9DCCaGdSiSgpB/EuxB1Y27jnXzaav4dUxKDxw1a60dr7NUIgK2Vztcl02ajf6
ka1hMkgQe2dnBG1g53XTR6Mx+tNN5Cmytq/OMQo2ChsPvpkyki1BWuXC0GQWZk4KNIb7Yqe40S2/
Vvqwan05T3ccNRl3/vnWW7n1t7GaWhfjKCEVXPaT6RYX7s+nSDPFhRYP78NqxUkKioBSpGhGDbph
n3ROks8jxU+NVjoJfbld36wUOBTqVyaZk/7/TTBKuT4jwiOljPg/v4n4XWFklJzcGQy4IlecF9tz
9Cvklbfp4+aC8r6YtSzKQhP/czu77wo1iaEqcOYMPO4nvdgDFfSibQ1OREsLSh13J0MCINeio1Kw
3WkXZ/0zS0kpJM+KIbVx2TfuASLfuNYjokz4LwvoiVamdUkIP0ygJkc+bQWmMbJ4MaAp/eawXu+B
RBNVgSpEG+F3uFOvByc0GUXgkujx4uR603xO6JTYdIq9qDkIgFEiye4UZZr23NI8iHmQcXlX/aTY
ey3pNfC6UcRVsLwEh72+PZ6ztaMaaZJnSAG1A5p9hogIjz/3xhwk8mxpkC3RdzgFtFWkTBbh5ltB
W9W6xLVdp9K+R+RF3/yLJiMxqh2D7F8pD9oc2V/UkjigqjhlHlqqJhLH4cn0QISgC1LGLfTrY2Q6
6Rt9A1vyrbdoJnf7jU3ipwQZXITtBQYGdOJWsCoTydq4bx3nQSyqZ72OnrESvMNU6NkpNY1qB5pu
PORCYqCWGxDH+jjKgfg5imdhM1UUuqsGWQpazVD7tnW5acuR2UFe1+IL8BaF/fVRpQmv717wJWeb
t/SMLV/jWDW7UuUaXcG4KUivCHfHrI0+wOCV0mQqcZRJJfhXbu19T6Y5bWV77lUVd972Er4Wv4Wa
/fNOAtQblg7gp5eR+lHdevPwpiCilhMO9SJWTJ0ojhl4BBhtPIHr6O/Lx9BgohjYJRE0wwVQl3l5
bFHBegDqSiAIarS60c99nXW0smCsYEobj3f+fcR7wZTwWLrkFccNh1T/h+vDayWKbkQrqf4ouMAy
8Cw5VBPDdT9dxgm3DHv4Rthw6IG0CrkQVyyrjPT3yPSKzDdTZ1p5qaC/d0y0WBlX3iVGwL7PEK65
nsGpKG9lfjhRh4czbTWg36VdnSNyPtHL7Y/xKO+4Oq8nHTd4ITOwO10SCdOR0JcqTsnh6Ddo9w7N
OPmbpaKW+g1Mhg0dcqdiQrtoFxvVR4atm8lNpYEKOCxHT8jLgWzfAu/HML9EHfOSAHmyRyMmMtjZ
BVZCW5GUMjDeEzR252qnLPQXfaw0A86GWkapA+G98h1GqUvKBcXWNIrObkgUWZgSkgAS5s32Seu2
ZaHb8KW3mfHVHQ+vgnBhhQvGLb1V26sB8MbBCc1ggOw6NoGWldgLknG8fqj1XinqTOCyW1g7KNyp
8KzWNKp5OCYV3ZSbKTI45VpXWnuNaiXeGMlsgW8vdPKQWJM038wH66MCiN1fyrRW7flMzE9fw+JX
n4wFTXwC2ry0HZOw3o75b+gMI4BW6YGiI9nC1nZoI2znrJwWvCsLbjelQNo5L3gB5XeaxqoB9d28
D7ObSestXu2Qu1A9YwyTt8UAJx6dI9MmYjEvTccCXIyvrzNOAWjapf2bhF5AhCrMXDOxGvhqdllJ
gYT568po4/wkEpEpay9+B0oFUeH9a9lWiGiROna5tcz93+t/OiE1KqWw4NCU4NJRJfdMIQSpJjuA
ABjyEqUlpqwirGa74EScyMAosyNAfvoTq9tZhJxb7pbjKD61pvoWNYbjMBS9xKAA5qJohqyiBcNu
M/j7CnGLT+A3IIxB8M1uWRu67NkALC7XY86Enjx2j+8HdtNEEM2QIlyPmuK8WhQeownLEnDv19Lu
Kt8f47qLGZMMx5MYlgQwqUG1+fT8Nsgk+5jOdtaVhAU3b061gJQpxncIhNLw9QQm8aVFe6phpHUL
2WXuKGdPlwOPst3qza8RTQ1zQ8hE2QNtXXZy9Z/DJH57thrysHh/9tyV9cVuhgNcoRULg1LsUom0
0MnN3Nsl9Truc/mmEUVrzRs3Cdx/JE+2cmTZlP06fVCKoj+zNzFffe1I3fymOF5PdbPVZHe/bjOy
lHi+mPSt424KoTK6xk1FHKQcEJKwrFYn5IYmIwQw3CFp6uhthaGCciq2GwCwQ6AewOQJz8THIJg8
MKA+/52+nCrpQ4UTZtzG/zJkI88r+VkU3IMPhJdrbnrW0/VWszbjMcQ8wvgemGEWQdMRwZdn0vjl
elgQj0Yk1ECyIH0ZFDbYmD+pJ/KI0id820P301gquEidXFkn/fkEAEp9r+mIzfa602SqII3FKcjI
xUARqieHq+ba8TdpkYPLBlRNBUTK9sDz2H6RIP9/IjgUI+JORwAlG6ZdxmMKEUVOo6Mk+ETTZIBy
lWjMB3JkbWNgEmuUMLHY3UrJjP5Qw1Sng1YySBH9Xb7iJs4Yo3GRd3lzmD9GwwLpm4+SiMeVu+ZA
D65kHXcKbd9R/7bb9+N5Rp7pbIL/J0QZSQXYl5eU64yxY3/2EEzUP2GwNiw2Zt6q5h3RYZv0AP+T
V22q0Ces6WEI3+7viCDXapUl9jD0RABe5/PErQ3swGgvnuxXRx/pT0FWuWS/7yTIsoXDIatRPdyb
RggWJiaYYQa9E+NQvsp2pMY4r9STwTEUeFxT7TidZW+guG8HbfKURi6HFN8suo8XSVhec4WO0GSv
zZVgfYLqU3ZAxV45C7b1jYrSWt9ZSC4Dh8irAtV6AIFIxIOso8V135NXVutLOGcYGziTT3crPGsV
v9sw3Q4BVyF/2uutHJUS4U6V6cvbKH+GTZxxlKzaP0B0aW55TlZZ+5Q+t3QX2ZiPku0St5e8i+Ih
YBil1T6SEW5jhsZ+vAiVb1aCySLzzSUgce3LPwnmOrzclfq5+WJzroOstY1hd5xc7e2oPLKnswvj
SLWDUYm5tARq/rOu6fQrbP78Dag2GnIWGhMsmdEGNaRIWYvKPsm3UwnYkC257jGhRgAoUVFdmQnk
zIdLQQkcnJbgibxyaIz8sVvpAhEDD2mHnkHT7fHRJvQEvedYocJ/c9cKyCRzozmic9jJvqy9vWZy
UYaQV30dGL38w3gaokGawNz5fidQNdII0fAjlZQbK3iEOCLFFEQFIVrDlJZh+squWV4AgA9+l/o1
PV/lBtPPcv7LZlieNnaXhSKXLjdYNazg1CKv4yNX+YoW45lhR9uR7k6zD4+UoKdtgTs2nQx4ldcr
13rzJ6oYquOCFnqMsCEHwNHW2Z3x3g0ei5hXEvjQErV21JNuKiJB5U2glJvoJYoJCVkAHLYthYNU
jXMwB39rYTB0xw06n0kGiDiPjGJnBzH7bx+VXerkgPX4NCpdehzeAKFq1nvubi1GSKXcfSNb6zNy
/xS45fgMVsh0Wz+Q148XjQRplo+EZ/AKwKBOAi7oavWtgAbFcdUyky5/2ZM50XU4+FwwTjHwGY1t
5G9Rt6e9yrDZFLrROXZZmukjFNUz4T+P3iybJt3PcmZW5Ee3clMXz9f3/maixQk0IP2D3/6b1Dfr
RaK+Y5ymZEL3NoOMBZf7rA/yQlNvQ7mUO6GZQPzQhTmu/rgtpphlR4KTx1DJgYELf6QoNZS36gjY
THWDB735rTXvVroaVDF5NaAZx0UN+La0BIKX/ik9N6RZwZfAJ5z6bpTgqGP5c1tqb3xtD6OUZMsb
095GHzxZc0AwvAtvpcdlMH1eqGcC25k4hxX1YDTsrilp7sUmE73KGh6c3M9i8rJm5WC7MTLp8JZ4
yNy7WZiZNYBN8ePRH7TXbBXI70FWAeSe0rJYNvFTC+xbr6NwEXdSEacfWf0Qd0JHNvHgnrUJ1fd1
uUnImFnpgENS3ltG/GMkzjXsEy04HK0PRUNbj+iWlRYhJydS7G7EeCGBuKp603uBwxZnKUUeqk4o
RQ5LdExBL2m/f63U3K1vp/I2cWOVlVgg9+iFAItpO0iqfQuawYjUXDGIFRNJCWvOqMj1fjnEOAQO
Ta0mVtTFHY2OR0N8RcQnDOxzUnzSJevEOivgCM8jfpLUeqQQiNklD3upBEk4iXs2QKD5DNUAM5AC
gIVgFBy0tfjffp9/oVtAyf7esE26bwDS0EotE6SlKst87J7jfKJs533v7cXzRjtSnoayucebbt10
aZoSMSk6J2mubyENyy1E5vN1L5bOY+IulFDjDIaszsqmdyfxlj9hmd0+n0rnl8rCi+Ecf4EP+Z1P
9nasATaafSpPxAGr2gvU4mm0F98tsoU2lIMiI7Rqn+OcT9eDErcnrOHrEDeruRztv/fc/ND7yqPo
oPyJqmv6rwKru/Jprx3Azp4wgk84apgri26tj6ny+5i/jTp9sgU1IOQIubyVmHGu3tlCPvYQFYNY
pvKi0niBbwzDlTLFOOh1oenxojwzODYYUI6wZjeXTGhv19AmdkdCbysrsDtlLRg07AVWX/7BMets
mY8l9QuWiDLDwMmcibw0yiD0IrNPxEEzOpXVbqkeLvXp3NmcPpu8TRc5OIxEp7M5WzI6FFBke/Ng
LmhFvD8zZq583hwBSax6JPxqKg2WRRi69jhJ6TCIQJgJ23YMqGJvk7/iWr3/ZtqRB7l9oaEevsko
8DM7Q8nfQ+FX0Wf+K/lYST4VIdtU/EFGD1vdlrX2NpmPWe2zIvTIsnhatO0uKnkWOXHncHD40f8C
JHFNfYLB6DSfcHp2ampRkgxfAELP80P/dA/eoEzkTAdPsATLFKUiILk+9P/Az881PZS0Uov1A/tv
9RaPcMS2Jd4dhXiH/Pu32sLeaHodPRpDwf/k6vB+17W8ilJRpYguUdjGP98bLzzNXlM+on1wnMqc
MpXAAqe6sV1841v/OJQ0VU3KfTIU8j+M6TvRiZOApZO2MLQv8kc/FkQP3lJPiTLcyfJzjEvnYhOK
Ndw6Y523kwWE/keUJdBtC9Js3CqtoSIr3weQcrL3hBzqsTyvY9s6MW1B0P8QQ2bPEd546iiXpNy4
HAD8sTapbgDWexQ6IbawngLl3Cmqdz2yyt5pGcO92XYTGQJOrpKegcF46G9TGfrqc19KldafNxcf
0BwmTS2L1ftqSyY1HvSUftb3WsbSvRQiK1MWOWOluOBTHz3aRZGPI0ibnnjGwOdNrE6g+qfY0GFD
66NErK2qaNBesSdPr8+unr/sh+0C6yWr4wNb/hfsnE3pcOdSdnu0uxN3w27fxs2+lwpLRzYNsgoA
AJKrphLh2oncG2PoDiFnwXaWoMSYYXEU5LFiCFiAcyVN/io90QtH4cCud9yX5Nu10Rk2FWny260p
UtyE6w1AYI2KCI/Ay0Hq736McLq+e/doC6iqvL4EaVGW+faa+h/JaqkItJG0+xjhTAbZgeBNWfFB
20Y7aTgYImsdb+88BevSw0t7Zr8CzM/SINkKyNRUBcaQcfuNXkbGvuOcvQNgUqoS6AbjjURkfXfc
gk6ypBPwFD3iAIM0LXJPBG8e/Pelrq40gccJSs1M6nG6+ERxZSl8C+O3AoW2fw80LqZHnT7qiQyT
b2FsC728GN9cKBK61xwNQAY31SglFJngaUDhPVE+ot1DEJCDl24Fx4uTwrOgG5XWTQn7DowsQ9ZG
i6S5kKz48NxMEEqAsU+oRfhAbONtsDee5YO3/mhm5PEaWKu5a+0QLTPMlTx+6TSMld/JS+meagX/
3JtaV/ibHOgNmRVbE5DARz35Vjq38Y/QMOK2NqoxI6qtZ50ufy35o/g7+eSUTuEfPl/sVitqSjXv
G6GFy2kXaAWzw2k5F2fLWvQ0BufIOH6eIY6MME8pBhZo20xEObQFcA9Ur3WbCHMDA9cOM4Giuyh2
Q8qo2DCVdo0D6x+OkjJ8UmRE+VQk+GupyuxNxXkwiKJuErDcjsuKSZMnrJKeO2zIlK4o69byj8tD
34zJ1/wRYYmjelFZQjzChLjKm9J/zVFAXusy0uFxhRDK0+4s3EW1Oot2v/ARiF0T66OQTXxivYZS
gP/pddy24s4Ck9MISg9jgdxmoIqjv7wzUa4sAlgysRV9K4lXjntpVnfKmp8B7EJew9L1OlrFGhhH
LCTsmbcEoDvdP0A6xrH/iuSzCr39TL4Q6kAFYskQMwxLM2tnaTMjyziqgsW5AvzoxAU75Wb6kxDc
alNqM7RWANsFn2ct89faRAqfFKEj+JuYwtbMWEh+johdyM7GcymCXyEEwLhDqUGLmVvvLheknSbv
/3xVU8yS7nWMka3GdhTeg6sj8XtftHIFszLgO8x4wGYOmxJfGeTwnOgDE7NfbxulUgFqMv8eSJCJ
Gybm1ZBfZh/JXLzQssFcAYfSaKSeV/4f6hyV57FBgZaxrP1O7flnHKMibrLsQcr4EhVlHpAk1hz9
NAfQHzTm5xCSIMNLj/UodqanbtiybBmV7XSwmFmbx+rDjrEmV1SrkL8QnWjS8FkG7n63P5pHvN+R
5PWSJEttxJSSjsbmUkMjFqQ4IsRqoc1QHaX3iSDC8wf3PENnOSWUnzxZ0E3JnQDyIouK69R7AViL
1+gf6F/jNpBg3FKtiGRChDV7nq4JZ/8layfREarYQ3+YMMnqwNdx5OeQl6eAZ6nM8E/OfTYekwJK
NTkp3+Fec9Aww42cQTCtWiZAP0Kc2MSWxlcZ6NSb7SI7rdHJopCxBxoBd411qiStukisy3OP8p9S
hEcNrwmHGSt1H2YmPdPHMowDIW6DVo69WMkjtPCNpG0kHJrsESTTuQEvXUt4OgTBkj7t0ws2f3Ih
YwRkgD3HG/RqL+WYrVB4vQ5nkVzdJbCIBtOJ+o8E+YjDDwVxgg1NPHXzJgyFfkO1khQtaWbwQjhH
kvSc+yBwwre0kg5WZ0IJLuibqvQsJ4A1AOlj/zkZZw/aqHy1Was3Hp1RkcZ1lkUMBZskO115xYl/
F2qkkd5+jcU16Ij5+g/CPYw/R4TiED8GV4+5PU106h9mJ0BUVp0BkSZJCggISJc2x/OTbkqOv2y3
y/N44fR/c55HjCllEnKAR8HS7ulocQ0mFVPadm0dt1zdjZ/ZEuUkmZhf/VnDGBUOpPinPBMOJsCr
nouYEKJp9VCUfav30E9ttKqRFMsYD0RXsUdToY0m0pBPcjTJ32AnuyI7iuW+XsC2RrnjnfWWzOyp
AczoCuKvqb03Y9W09BamXtqTm/5nqRQ6d46JYteCamvAiOJV5GGIvqml8MG8ORw14IbG3WhWYW+D
IBfJtyT4Qqvl3ckb2WRUk4vHRwrM2GycLG9mseei5T40iJNCkCnnzNvI5DQmUDQmgT9bb+pUawV2
dZr3Xy8ORyomqbXU8w3lFnTRsC9sMDb+YuHXZSR6UkvYBb4lQxxyI6oPxnEE72H2e73pgV4jbDjo
+879qv+XVbXYAHyBAWs4K450mbZm63SSC1SXNfNrv07e1ekggRjCqYlzFnWsFC56x1H3c16kPojI
nLDyYrygDxTGO3FpoQRDHPNl4w8SFutU5cUdeL+ZvxrokXfZ8BVGety4vngXVFXPX0xNzFdeoMD8
2PnoYuegJaRO5tFnfZLnv1R7+5huy1bIHxdZtZ0OW/lQev5ok3/ebG6HiWdYLjrEhWaUgl06LDYA
oxUrlwhZAPrXdZ2EGHP9VYZT2O1GpvzS4NEO3EY4NunaypikDpYmNKgUOcjHbmcPy+nO0pNaACGn
LXeIgLTHrjTj3LvyIf1KjY3/fHQ5DGYeTCbkX/g+tlnt94SwhsLZO6cegkROlswhNHcq+W+mS8R+
cGPREzErHB9jArRTvUTfscZ32VGI1yP/VII0gq7jEKflxomRQneq5l9zNXfBsxZanOAxD2YbBn+U
0ez3CO3uWs/fckGkfO4AeldbEDlyeq8Tw1tzNM+qFlHhWIrG9iVInZN5/ydnz7AiDZonQfVcvZ0w
xew/ul0hX5x7YZTOZ86eFaUux5MTZTMOUGxMDj6fxv+YVg39sGYq20wuO8gVqjLGjmeyE0m0DVkh
QlPwcZSjlulDJwoFP7qVlnwF16GOEU0WEoUZbNaY8sdWjQ/JUmtf36ybxCLX5x+hX0rKI4Bga70x
H28Eis7/N91sNVV7qJYim5Sku5ZX95WxCSd/Vmq9kaPmuRs/YxSamDiLWWK8p9u24+HLS4zjaH95
vdDYox2Zug7nvtG6n9mx/T4/em9eL9mT1xuazvfGE4fLTSok5KarCTQspSJWazUAeHUbLzIsQyCz
gWQOB1RR06QsDXFRLOn8tQOXYDBcrkma5QSb1h9l8ooLVeHwJodtkGUs0/4Z8QIQA9k2NS04GNno
FM8EXuai+N2hzwsz32Pdoqyzy+5Q41bf9KWJhc1M8eqeLY09FHQ3WgM7DMP/kxDt3HkSJd5RITB/
vHFp2uhmbGGeRr6NuieQtaiKYNuJ2kKLXqVB0iKsDYZi4mIdyKJSrbAtvQiNOkZF6RtCfluZfn8S
noHEmqNS8ZCkGvI61Ui3EGjQ8rX8IAE8Lh0hRBDOzx8Ewky4/mmAAa0By8QaSGxdu/j9rKElJduM
OgJHJCj9IWmPY73+NL5q20x44Ve4mnuu0OYcWFy2R8dqm8l56kYiyu/tNwkD4LN3QNx/gQVsQm8c
6B+Vn6HVbNp1KqYsMKfQBA33UIjwPt3GotVhIcZUv6Nbh1A9H9FV3iEod3CqaneIR6WhmA/9SdQt
AdHnvg99n2nSDutmm5g/tL6VXvordzEieEmCJPR/tNWNmjcZA+lH6qQynSVoNg8vAMgu1zmf51YD
TtNVd3LGYg0f9Je3kSw6T7FvOIhPgQ7ECT1Mll8qtEUbPXlQUXX6iJYMUMh/ITwVgFd1XqiiMQWJ
7WNj+/ZmxdysGiy6IZNtzvjiEgyEewfmUA/PlWSqNRfwc9KKsCqV9EW1hNcxQpw8rqSOuPjFJtpB
XmbYtMo1H/MuZXB8VVTm12ZGHc42SmFGTaI8UiIkhgard6ujJw+OLuMMDUMLk7mlSNZjkjLLuIaj
Zzqu9hrloLtzzN27nC6RPfW/OdT2brKxskWpIdK+JjkXSSZu1308TR+baZvF+LQ8R6PAhXI5uhZ1
rexnDy4sr8FHE1kiiE0uEYDbC6CGqpv2Bjzb1xN13Da1EY1JhAqISzv31sFKhKtyMXnUs4pWNXDO
bx13YCXEgQ/vUmWtvn3OTKx54kjCkCF2sc6TSCXsMISpYfhLxwl6C6csjXB0kdtZZNBnF1a93PQX
+/BaD6ONg709vQSCp6mYYih2m+aRubr6hb3iH1kJrTReWMOXdcJ5KNzkm/PAd+p3IrDeR1b+24TN
gFvWWSfc1RqU9LT2uLvrb3P4AFgQRL8mGvy3kE2C4WmcYCDtpYOsk0Mdc2io72ldZzW58/Mxdqvr
IFitIZ+qmQ/PqG7MLezULtipZa3YM+8+w7VppOap5xL4qpVO4aVUoPFkIXWk5lo+vHkPJj/aUz4j
OQ+7PnV1lEhv5MWwy1GAna33qua2dnLHBSMTTwTIA/g7zfIuwbUn+5ipyW2BvPA53GnKYTORQyB9
zkYmAGkCXNAsPhL434QfOxi0GjskARPGZZtBcxp0vsL7Q8Wq1tHVm2sfX4oRrPCxjfewjjudNBaa
cikScykFybZ61V3BeeldjyB+yedg7kkFWTqVWopal4gQ2PgTqeyFMIZkactbtS1BCaSJpyosD3CI
iwRR257xJ5B3IAsc920blUd8CTNjBzDckiQ1bHvnife1YJNl+BTNT5YFYhoFJqPKwi2+vGXCIm9z
o334WHpfFfVCiwC36+jJHF7dNgvFHCBjjBHDyprSt3fV92wiX7yChQeUz4OkF1LFZ9vKfIQlUiOy
UVHFiEsWIaLk0UVFqpe/sMoetx7+9EuxtkBgjoQ2a0TnaJUydFpO8dYH1O6aPlwWuaod1/VNqd5P
AXV4ovZaYbuVvh1bJXkO8aFhjhwfKt/4yWJc1tr6UXh1uMgA3m7KP11UDTwm1bgmffd0e8tSDA2r
oyaSer8D/JyIVLAy9ePoGL6DSD00eUtTz7+8MYAFV5J8XzITb6rN584QBFWoxyk/Jv395XF6mDv3
o5Qb8uTZNRTRd6sgZJJ2jocFMp9AhiOyyv4YndAvg9jr05Q5NGiRH+DU3tPRKvRJyFwpyjvTAZTl
5aC3u4iSmzuV/QBEV001ICb2Cy6gFWO2rFYo9ETzLbGJoP+QqHVHO0gcPKDHn/+eQIG7b87jV8YH
YQDhbQfmsCYLUm3JfAVtnyQp11iG5y6kTLnDpmJfgBDouzGXN5J5TEGLIqxLZATBYX4k0KBtth5Z
axWk/lowAy0RmNMMlr1kW0pCmzMc7ZByii2EskwWcJXAEiGB7ZbUOBcYg6XPxKMVGCcSHwR+xRsH
QRGBcaTli8ulNAsBgp83o2/NWOEOs2VAJvolVU/kBg/AsGrsA5SxzF3ysty89DqJebIqeZbhd09y
a3xjnWqf+cvajh7Nura//2WHzUvhK2Zg1qJM+SARRm3PVZn98J2VDUVj5C0fHGGau4xuXltdhqSW
CGk2k2ajHzrqe/ytDNdeMXRFFi5IT0E/In6R5jFsBti4m5PrfuSugYEx+NMcOcOzN7Bu7qn8f7vD
wrxIGep1vmQHJk+xlm0rCDYDOzAvbX5+0ROmMtvtFLGuypsMi2/Ja4LThXzAyoktZ6Vq7m4HDhIa
Ps1Nt4ZmcPrUjoao6QNVXCxFn4tjw+6NnVqEp9/7lauWPFBk/wh+A6yaDG6teSmk39g52lHvLxpy
ZWQN7yQS2YW//LtWWWeDQXeiVHqvYnzuh82jipRtDCEiUxUCrnrA6iOhOodvl9K4zaRnOoTry/Yh
V2mcZ43TSvuQlLxuKUDQTGAyvgWKLdDmu4+7YnEcKC65MnYn+fSaqH/NY31cN2lPbOWy5k7KeC1D
xa/q4lHRo+gx4SuBiy9bPJmomfNw379/BWlaHUerJJZK1UV4xXUVTwgOAFxrxsuIJWxadDnAIynQ
q6px5Oru5/4jkLpLHNO+A5q3x4MCuEQoI2gbc0aZU2aUNny1IUiDU7G9d0uYEx9F6ojmBj2slZjL
3puqoiVfqEn8YTCgOsp9TGsHKS0a9bkVZ1m8wc1HUn0jO05bkvxhg4dXUg3xPyTXZY7Xm2z8Imz4
uRoZnN92DOmvPHaUEPlxveErlqbroz7oIKfMZgE+1iTWqMYT1LozI0dpJq8FEvk+65MgKCyhSbJ2
pcZ5YsonU1FjCw/Kt+Qjwn73rRs5e+qIS8GhG74NBY41wXLaTMcQ9ZW9jYduJOzRX7tCfi38xKoB
E5Ye1+TyY6elV+1KF4WOI65/cErwL4RLpde1W1J1GD9AQrWtGMhN0iX1vD0wtLx9T2ZVt07gPOqV
YwMLbCEBUQezt/4sLBFSAtBkLREyo9mVd41MonIuvvqmHw2hLfPwlgVq1s46T8etq0ab/aRSEKp0
MIPrLTpvRFckNj0YUJxwC3IOqPXJsMpnAcallTDuYPxtuS8iIkRJqq/AJMrhiVfoD0LibVth2jDF
pWr++CncT4/kW44ktB8i+VkmO4Lancj5Z1NOpmqNv7ApoRVoXohWPSVWpjzeCwqpTiyo2RQXUK87
Fnp5Fa03/OGcoq9y1JFQXRhdSvInG5fVEPukPjOQ9S2s3CutbWrMtWvuTeMDfnIz/aZJzgQIcVXU
ySmXA/L4RkZ2OFIs0cVifemBw73rw0WC3Z5ZVfTh8zN1d/zAr0CDPYg823KEAqiTQyDJJW6T7OhU
hzmJfwXjLd+0jIF3+ZNWSCmM2v5i7fzoQhz5j7GrUxSVRyFzhKEUzdRFkL9fgrv92Da8vBZJbBXd
wjfUKWyqhA2mzra0ZXYQXZPydoeHyd+MjvXDuqkH0gkbg7b0iPgLInL0Qaz+6fStFc2WozZ6t0kp
9up9ApTkMS8c8QSom3g9dw1x/hfTRrIA9RYfv2yl1ZV5V2O7ur7AmMbEy4vVHYmcDcRCdVcj8grM
1B1WjrBOwQlTNNzb9NHsPrOTxK9LoU+6qkLVIqEMAdda4Iqse3IB5CYOSHsHfj7jqPzuD3AJtU0z
qKTxnpk/CtIolx3BnXZ7E16FQSTVlF18ZS2fQaubvD9WnTfW5+AIgtlXhBzYYAdiQPn/sgHDNoLG
NOXjDrANtrfUKV55c41gIEiTVJdhG5EmKJlMDkRBP8yjZdQH7tNPNLfCUEch6jUHBd4Uyv9Uj3a5
roK3h3jtn5IdHkaQ34xuYfX+cyI0Qn71uTutFzUSylkJ7Fb8AdLzzQXonrfetmePuCObyzxT6emh
nIueAiP1k/dsx4vTiMcLSqCLzU5/yMzgICcHzzNYN6zs2wSOJxCqLL4ubseg7h/nRrXN3ULMpRdN
0Sxst/uAfbNroCBdLpDbOBxXCI3yOvkIzdWifHV9toi2NcnzY55kOyx0GdO+XeCu6AewBRbuwp+Z
xoEdvb0cWUFFbQi0k/Bp7KsBW0AUfGt7qjiDqPNjYqutJv0iQMfgbW7jvug+O0kyRsW7Rbs6yJw2
FqyLkla7i5ZwYoFsQnArClb8zmnHg+pj8ZV1krsxkVVjO0qxzwcouJQt25gglotk96B6F050hlye
kRZxM+5rl3eNRoXS/qhltCNxCR1qH3vA3KWeYuP9ZzlmPkKfNpq+2odphd9SWEIFYlpfdX/sD+Vb
89nJqDfUgwO2BOG4/D0IVSzrqO5hsYizIWbB7M9t6N+4+hmB44Dde7Jk6qOrRP16mKyLpGyGO8xV
5+prIgocftTocwAs0Oa1Hi2TEWcbLxAIgivQo6Oj24l6rJvbInBuFHmfZ/cpARGY+sO/LfV0z6h5
l+Y5x4en3tQeU5vIcW366moWTOzSUAzGaO4BLRVhGhV9E2dXODOiQvnvo19OuO7Og4K0A1LTy36Y
Eip0WG13w5LJ2X2PP5Ila1G2lmKGrMAUEx3/vgt4YG7x9lnobvpUZwEhF7gJy/Y+PL3fkqh+LvXb
m83IRlL9jhnxdwojGVAYYCeg+oIcB2OZLRQs8VOWJc3hN6g8DEW4br9iOSrQuPhT4hFPMRgaZdv6
fx8261fEkR/i75erHiBzyyZr+bFRHICAgr7FGPNgt4lIHrYdDgO8cLcP7NIBcguetdZ5XfG9Ae3a
z6XkmgfYcFt5i04Xw24acxDSF7t6pT4yFAOGAJ8kpIpEhR29WaXTypOdShPT7y4F+RdpePJzarxx
B4ZHtfMU0r8kFt6Qsyaka/Mgud5rBxTpSrrG5lqaZ9iBH9LwKgSA5KWgEldbIjB+nysiuu/BZUTp
//NhOixT4WndDrJ+NyV9H2LUzWfGvkI1NSrOEoMVttjFHFVAM9JlQ+G36h72gVVGQB/nU7FMAJug
7ilNrOUvdFQMvgIf4lCBr1CbGUKfawQ06NHvULjcu6w2GaDmCXpzUocomhDmDY/0/O1zbTGJ0iGo
xDlXTlXAnZyL8MGCTGBEC6UeyNSytaH0/gZIWRhdTIzgSKDR3jfysIKGyOVue/Ei13V9tKpeISuj
t/a5Nz7TLtan3lyBMxXHwsXgVFW8z843pxtCOwaX3IiGuMOtQOzr17++6duDrmxut6QUTdnhS6Js
kpRGZgUc28rMhoO+DSWZU00R8fgvW7DQj5uF5AVire9QmI8NhHCSkOULhvP1iUQMkEWVq8lHMpTW
rpEOEQ4uKM+ulMOa4fCzmyWdFAyAB0A8gEkhoLJgnnAFaCJmVjU7YSPsnH9wxYx2AHHeqPXYt2xm
aCgJzxWqady6kzAQIX4biHY4L7wj4EsQaOhfWZf4YULL/WEK9K/6Z9dtJtGJTnF+fmvEEr06+JEo
EIJBKXKdUDJ1h0jP8g4XAzBItRpD4ONhxAEltt0hoKPTeR/mPcjJ/Sv9cFKkuePZDDiB73U51rNO
/yT4pfXZacM7okJwXD7+YQA5rSP2zG5U56lZCYB+tdUdGC5U4pBqsLSPdFyzuIV3JoBos5Lpm5HT
SxTVjQFOxOIH6e8Unh07UiLhhfAKrJ8Jx0JqPkiy68UyWqb3ETTZmWr95XvHg0bWkazpyszdeaAe
yxfjoqM/J8PU1X+GoNNhUMyGR4e7iRl4wRscG3WUlAmrqXoSm0BzzjBV3Ie6RVJNiAcjYh32JuVE
tXME/PdrXDED8klwPbCa7dnw9S3uT67LkLS3VP1NITCcr96YApVsOirAiTi3h1heVATQ/aASydOo
cjAE5YzYJuljJTzDMjKSjlYLVDrQZbdtYHRqiX3vwXFBG21YFHmMEPF3oN1AChMcHB/hDbqRViFw
o616AqEq3oC6fRONtXGynSHRKsWlZEHArWRZmbyfmnXM12NzDRNLpnR0AZv9IGmpZNTlL9VCtxA8
HPu7bxKwVhc/32+LlA3FYEnepWcEOrFFoVpj0+Dzg72PsDPDgR0VwOhalU9PZWHztv6fStLYrXdQ
bW++Bk6kOIJoOVkdCj0Tn0K5Dky2OVEjlcfPsm8E/ErDa8cz1+zQBqWehJ+UqFfdCOxE1CGLZXgg
oOVB4KLUqvUGwWKw+UMpLHStlrlKi7673PnswYXKvgK3adMblLLuqtWUFSKidbGPGM4RzTkvdHH7
5Nc/r7VpZ1tzGGaEzEUnb5MsJ5jx6TBW/Vcpm5g1k/5CgJ7Ts1lRFao3kCs6YItgHt9I+FzCEd4G
HcjparsTZK+0q3kqqFfliyLFmTAgqbgSixhJxuaBJb3W7TCVCutl3F+eCnnY1q86QiJCM0q8aanh
NTOAjOYOW7iWyqsapFxg3cPZMFHF2ekfKfJdYUWc4geguCP2OuWjuNdIYYTZ10AC2hu5kUGC6bQ5
4SOphPNxDnFmC2AjEoWVDw7iqGWPCU34Pvl3/n/SdPOkXAc73vyjGn1OQHXQvyrFWsneLpI74wkH
IfbQVmLQ7ikudaySDpnyHhRAmBFI4txZVngt/itnbO4KG5Af9ireo0aQY2EZM5qBaapbO+AyAjLa
ezEu7TSVTJsusc4XifVM5EeOejJ4WbZ9H4Mo1b6iHOLYxHKkHFUfKXIjnV38pzJ1lJm3rEa+R/B2
mXi0fyEq3YwIJyykIejVqBu3Wpn4y7N7JVKmJYll90cl0JBnz4j48+31kMmlkR1bJbIyNYE1w1jP
H6XS3AjkGOXp1oBy/08NJAmLh2miUJWzIPxU0DCUYa/7U7Tsx8JKsTJPZcRsIiuefhisatYT3EHb
b/wb9uixKry6v7PgE8UxnONlq7NL3LbLrmqEhA3SESO0bnDxZ1Iv0n/uWKM98riIPbkhQi8V6d07
vkLevsaJxC20o4bziGTzXyWBxzrnGeJDe8WUW7chNLWprxJOUarNvZICVrq9+SyWWsAj1kjWSCgf
2dWWESXYpCV2/w+u+4PxBwDjvyw+u61yDTowtHslJinQAok6EcExHS7SxmLcnpLSj87hk1Us2Iy0
roZjmpjKKF8ct0tm5+ucbQyqNFCZxWz2EARcEnENzHENIT+CxgnyP+a6MJMdMcufihJRYjVDuvjF
wniutCASzNxIwYgVdVTp7Xm4UzWXbhsbqxDwS20YVq2AeQfCE6muKfHlF9OPnSI5Bq/PB9XSoypu
QcHkXn4yxR2ExZxDkNjKYf3Qft+wRn/jbS9pIrEEVdj3lsrQ/w/vtQBqIw+PDMVsyr9bRBFJjx0F
BNPJAcrsw605Jxw+B1Ofm4s5W4hkn2xFmChCwDSt/NsSf97+BVe8y/wpfd3JXBAGNQBLiGQgkuSZ
MftiM3X/zmQ+1HtDek8z3nBOzI/sCPk/XthkpQjNMr0fazZaZukbP/uk4+ltQnJi7SFWcf8JhFxK
VciW26o+vLaTWI0rYAfXC3OawOKVoXjw7ePEkNhemtuDGb7kva6pxAmqVnEtjOCAvosejdMO3JJM
jSCl/fbEUvMVNR1f+clXbxEE9a13dexIlro5j+ODEZjcLCY/imyIZF/Iy99jvh7axaip6j/1Ah5S
09KIQImGaa/slAZbr4kMNhEcboZr76+5VyYNnrVUts2pqm2wwGFVXMzJkgleDiR+gSuY6mEZSkdm
io+8ioLD5H+vXsewCl8Mg4H+ubpEKzOXLUa759nfv3GaPRmAUeyAWoSgYEzBEwZlATbZVe0o3o7q
XAPePDbRpfj9Imp+dSETDpTZ7/xdK7AvC7rRbmqHJD9r1UNu4TgwQ5MJqcAcHi0saOMNSVWVNY2z
I/J9bwLm7VBNDL9qKxCNopN3g6s1AT6//dfFroy/p70UZDeVP+cf4PumXKWmsBXObfQiLdzZt2za
aGvDlnojrTBJkuwPBhEXhcLhgp+C4InHERLtRoMMTal4vy657Dx3A8VoUcB8z9QPj1EryDAZ0Iok
VRkNGB1de3gtuXzOLgQ+v/BfwRYURaqESRdGfmjy0VZDayJi6nnD0tifaXWLQzi4xPRNgqpM1b0a
2BtEWAGismdSbk9ZrNgdCbDpsL26mTmU/PjkLZpdO66eZn8cqUuclXIP9QH+dkgQ9OBbpJSMCQkv
mhqiuhf8IcP5CYWGHK0iTO9SnJLGh5NbbhKvxYPyuOeHca9CpmUC1zV5BTe7wN8g71yMrxf2HW/x
S7xNY3ccnWXBuBkGn2Uzq0blqwZE6jSEmWawpHyx0CE372mnkszvrBjXMmY9k5B+FgDy4E5phqOv
Yi0rW951NyhZSXFR5QbomyEAReknH4thsLH9sbrpEkqYZlccmv60NS6CS4+BR+S1mSzrd9PynySm
+nZzHKpGznbr+dDjfVxJMQXpSadd0TigTBS148sz2sgiPkR8XsEQCTn3NmAYsT+z8xeAYHqYFV8k
7dui5uMw46G3NrVRU88f4A7BTf4zQS1s3eNZsXgi0/bnvD2DEZbU2IXn9n4dU70MFwcW3OlJIwoR
gr1+2mmq8oF9abeFTBp2wk9uj6JsaNP+bW+f0eaShGXCY0splDcYwvKx9O61yB480qrFZ4OgAAj+
6BdLMWqXpyVmkIAMife2aFeCmkTURNU2wmSY8WXTuqKwNo+UGtFZcLpqtaJ19vf3LpCOa4EM/p95
8wUNbZD1e21k2We/dWvEJqZugkyi6/Rx1COQIAxdfeXS8BjcEgGvNydEWGDMxw22NnU7ruXyPddr
CWGL5ZPOweRGB0Jzpi/zkEJywl4swkQ1S1/8jnzh7ok4K3AdeiLTSP5g3RwreTyHHIuFY+OAyZOO
0SnIVl6g2uSR5iw9+bcPi3Zv+J2l0rxXgT2qA/tNma9DRVmgbE/9YbQfjEEuXHGVu+/ASLJ5BmLR
bMlSWK7dLAYQRACkf1I1NYsTyDBOw4Espwx/J+Mq5LqHli2j+H7TOn4TyijiYhA05PE3e1yymv9N
3M3VPLNtc6kWPtgI+H5E+q/WpqGBrnmSJU61ClwHDM2eCKt9Q9fgtJF3/KLL9OrdAfkkInh0wQpU
S2gCMGuTJKufv9Bo6ABmMa8zWfUzpKmsBy1cc69CRVV2rRUmi8Ik4PMWAOaqJahJ8Wq6JVbLxY+Q
j2oVpLROk1dT9TOLqAhUCppkrq5XeaAjGmHCD8AOgoddgEvHfE8CiBnP5/n8VdaLoa+Y48gIwWZX
54hZM1KG/T1vTowO4CPO7dNQmf+JB6F8JrcyiA5U48Pb09FWLUH+jpD0WX+BRl8vSLL8hz476ahI
thtDhWOjizh1Z+D+Oa3kcZa3e0ux+fxYJ4aWSw7+7QF2nxHwASYz2cClhVtqNfyeQULZpoiD9VzV
+8ZMqiWkjt7+mquQAgLiL3XJyEv4pme/ZVeVW57hykmnp3p+ljgebyF19/ZPRMsbviu3xI4gWsmu
uK9Oy24wUyncw4CF5q8M25tRjANMaH5LRdVWsx5i8yD6HmR3i7OtvLmNprnNCNGrHpMeQCB+LYtO
2ga7QWByLdcq6m1A49ykcWHrSbAqOsAc+SNIPzSZJMGqc7XgN9gy3lBHlAk8razAsMkuEEHGHc+y
+cGipD7WejWxjYBEG0yIi2ACZPagTGVO1yTLmHC91IVxhEw+BZNmhKpdRWhhyLhal2KNPFnBFylz
e6jLhNzhnZujQc1HIr1Kmw9WtzLwWpourjSnngmCHMIAhChI6RrjMyctwpw5qDiEL4cuL3TFEmMs
ETK7BQabw3cpP9yj8ZwwkGMqvgKPi5YG6seRZbznv4HeHHeGe4uGfuarXxbFQwAT6fknroo/8SVe
MrktKsw0he9gavuNvMvHBm2lvjQFgDQu7LCozs0bX0se/0kh756/tXvlMYy+qT4t8jcJ2jodGhST
aWx6QYtaucowN8aVUp3xMqsS/3BSHRb11GDcSvAWPeLXdktlPD2ondDgA0VyRlw9jJggj4Ff0K8G
bQwAFaDUsw2apx5CFWV6H5ekALE77Jly3A1DdJyVJSyWjZsjI9QS93VwD1/8/DCpJ4bn/zNe3Jrz
SxDBICkPIxwrUwLO7NkhTLKj/9Kx/2Rd4u7mUzZorCMGvn9iq9Zr33pPAmIoxm7h9bSVmKugEsEl
V05+Jl6M07MlwP6AXIKeyp21WdAMO9iDnMM0DLT7WyWofY51NKmVinB7usbVLGW9vo+mJK8aHqqr
JDC3RfSTb5KSJ6ZOdo5mXe/yLwCk5nCUY3miVh3JvaVAnn2OMnLlNyFi/u3O5fVo2u/+YSHmEchC
22A4BrmT73Of/H4wicn81Y6ki1mRSdPeEKXAhbsTZFunv/RKUNwP9EHCMnVLKDVpPG2Bg2ELlDFY
rLERBShfySDycZ378ZA6CeVs8gOMcHQMjXLQoBQMf4/sDYrPGJKMRaskhQDY/niYh6M5xqr4nQMp
X5ml70s1H7fpLWpUy5WlXBMwSD1hWOsIEiOOT/vwXsbjf5GPgcgwe+9rSMu53IYau5LQCTF/vQJw
d6UsoLnVZ78Ejb/w5uDi63tnmAb2Opm70lVjdtr3giPYNWdMrE6cM3oZYwjIal5Wkm5QHR2E0wh9
cp4+PONeF+MGmm+8Tmm0PFY4v+mQCt+ymyzxKVSBZ1lSb1jNApgxrJEFPdKvQ2lR7XAVwiX4qX0c
sS5Hhl29G7i9AqhFf7d9qYtPGq6RsN5AOqg96YNaCpfZnf1sEAU1DknWzYtTywxRfX5+/xMzVBz7
SKbmxrcu60LFCO8eeU03X4hz4+y3JWUnSK014Cm7n415HSL1Qw1D21M4+9yNkBdTnMmlb+3pYs70
tEzs3aWUQbnLscN0Jq402SwGIFdBln/h1BTGOaQYfxPv9nfJiZQIUVF6GXajWGv/p2aVci5jFfln
LkUCHo5dmReA25pL22vCfj2fH9Q4qPgY9WABDzz+B0mIdB5Qbg0EHmNbOAU0OQ9yPERQe9BwMYB2
7IfMV6ZNrU/Y4AtYT+RFoMYKLgWQ+yuiDsAD3O3bPWn1euhBLYD3sw3o3hBlnqlEeIL9B+TtbRgi
PmVywomE73/FDKi2OoJC+UvzaBM/UOYVVZx2B0QYswFfeVsrdR5ZK5q5sSB9gSJ+cxXpSQkTHTLD
PUVPKBMQua6MT1zAgXh5ScfJJxh8Vx1Ze7DqZTjcDU02GHYZiNhZkzwMsU/pYBCopu48yTwn4pkt
Gl0tneS1gYKBKveSflIP3TujrrpXqsw/i13E/tWTMh85qX11J0dypAqSyG+9qJhEOoqKq/E8wV7a
2MbrFoEI6yULsBdZqvgray1DRaWRPrbPk7sxtVHtGsCMaoTxFPCpyVyaRIY517qO7qpTWnnNpFPV
hNO9CZZvYEu2YBzhYQ7gdKEJMr9YUFayXIu6JUX84seuSeJSXCQssyeKhU9XdOLweCLyTLzMbn4T
IDbInFzI2R48vNPxMAtZ2LySHYrndzhmSkun8HkwOIn/eyBICX4GKINkaDYkdVDIC5WwDeK73F4B
Pf1h2u3herCZgbCBm5zAAhdODgZGgLncCEXLh8wX402Y1eo66oFdextJrkqx5AHd9qajsIyJw+mB
Tl5GXYVcRvdJIVHQy5fMTv5OBzxDeunQnV5VZV9SVnpIqM/tNwA9frnTz1C2RJ26v2dNrRimsgzn
gOVsaZdd+I0MmDtj9rSA7l7CDWdTn8k6A8pCBixgt9uUV7M+0h6EnFWgG2dRcQ7kSQdMZePZcz6t
owjRRw9pjSrRKH+fH0cHKnoj6SH5OTnv0PVjld7MT3vzGHQ2OUK3EWzip5RY2DbrkTZIhBOfYuvt
J48Z3aSwybWwCUS/Wx6737xnFQn1p8yH15tGeIlN5ybcLoqODDris+2k2GUZ0gIT+498mNfwMNbv
xJDbXiQxXq20az0SepM+pXrAsRae4jWQWdITXi5+h214lAcPUJJgxBHT0sMjDD5ySnRJJK6IOOE+
VKmnW5KHpnCmFMfUw9hXeh7LZVMVPwhmG2LbTaTw3BQO/l+wXxqPqhv045iAABmeDa/OLr2g7PSv
EptRLeqXv5voXpkibca8XSwulBHlEKLb+s+imBM1QNIG0GBnr9jkCDzt1LSEd1+71Zz58XgN+qVk
odoksO+Wg+HQnI7LrVaXP38/IyfXmX6L5WjxCKUlG58bOg6cEn/v2UtizOSvx35tvQcny1FmokuA
7fXVDihs0484BYt5hM5v+lsdGqSshrpOwEkwMMmMdamtza3+o7LVTPaABrXnH7A+xPnJtpuxyPAz
RarVtu+KZDF9otRzjG9wAj77PVqUSFPkgaeDIDAQ03DmdAH7sfWEa4m3JADD2rFlwU/NNxrUQlQm
ILcMkxkyoyNZynf2bIoo2JYNHTGaPDp40wv+xNyutNscgL8VWjtaR0r17fFXI2jnY3+8tMQQszXk
/isRS06HRpoboctnE/KuR2yUctLg3NABKJ1NYXt2KQYlCiOi8RDvRBzTnBr6QIBoQOvUbKgm9rSi
NFV4F8gzSkRIwOBzgB2RocSUQQPcfgXaEezXtB4yLYYZBaLG8oAgkx+rDFtTedMnVS/dZXNDc3vV
dQ2LvmnacA9I9vsFnB5Bh0fHOK3p5jXyjHF4Q9wLssp+G1HJUKZmGffH793/X/8MvuwjXPgliRb2
XbnxjLiTY3S/gOyH0sETc+4eC8U9QzCneHpTmDwLBTKpAzd0oHS84Ne4f/swc/DsUE1zz2NS6eab
r6HN1ctIEFLQ79FgVQk0OhV3gRXIFDMhUmrdfXvR+RPlgG6sewTjZiSICVwDt8eVKh9PLFe2QOqo
pc41pHQOd+PGkHnRYBIMdgFK04wMe8b2qpoImr7nvrQ4FjREB9ODptoPlFBNL6UFeNYWSH/t3GP5
EW7WZTWXoTRp34IgFns3kWu0wE0kbPw/XqjEzfaeNCADYyOol/WgNrET6s8dA1D46nUu22ya6Ass
LzoPhRV5Y7eAYiizFmDKsDofg7hfEa7WEVMHtlJh0EtEnkHTDGgg4/hi1PoDQ4UYmvLp4w0Gnruc
oHq2hVLQ0Tq9oAF0IfGLllP+kOWwzCFSA0zkpNGjpcdJMoRIH63xR1jCzkfcAD3aZgxqGkN/vrOh
borXnyYLsaszgiqZksj/NbLAmoCFSHko0ZG1kv/eKp/4f3l1TapRp2snqplSvfXzjAnAoDapsZPU
U7j0UB9/34uuzVGxhzplm4GsTv/MRUkOMLo75JEc8ZrCGAlr3PZOuxzHPQ8tIsedqDm2O3D9G1Yf
N0pgZUXhP9envhYx5Y00e7yN838IS/EIEntU/SzWOE6+MQi8hk7itmVaxXb6IyOZhFnvbFTVWUvK
V5lKvJJhSJCUr03U1qFHBEixLXuTFADo7XcAUbD1IP57ICE/tZKuvvHd+0IgBw8hECTwq5IsGqq4
90t6EMgsU++odzoiPTnbx39lG58sYzZx8BHZ3N6wbT+ai9sVSBMPe6wAKnhjDagE+u1zsvaIA25x
Yio0GEOMlaoK3/7MxY9AhdEqKrE3+hwZBOURiqOBm/m5eZh5rha0WpcnJtBUscls5a3ILgMrOLYE
wMnq4aXZfp/CQf0BN/3Iiq4N8latTTgCFlnw5YhhwKravLVgxYxEXFfGmEoANO5QnIhe84/rpsWX
95BSYsi6nj1SdM94pu9IQlBq3VHoOQ7Sb5MKh7cew5zE4gTA8GF0zGjzEMDtL8SbUAh32mBw+zRW
tylor3MX9Qkl7YbXrzyVzBhBFdm94pUMvNCrGB82ae28T3Gfzv3QoEM0eQoKvqclLcUX9QL88wdk
yOPVLezZC4H+HiDhqJsH7A1Z7o4xW0/TpIR+NayMMmm1xMCd2ItaJe6ua9I+ZdUHly1iiWgNUV2b
6q14O3krvkpl37zKDFnsatVLIGtpe1mKaq7NIeTTHD8OVzSHirsvMEVWTdKhTqTNDvzQrM4YRcfE
PWVTlv1jZxQojyp9GcHquxVK7vUT1tO90EfqXasTg5YEm7rbt2fLih1Kl/1yL0ubveH1kYweL8Pq
45jpYFPCvm03X/cTd2Vww6hSs5SSUaX+WjoTTAier5r3ij9/HL9sn6k5bE6J+EsSGkigTz3zjHkM
TvpuTqEqujvTADQG71afMuJWqn5DS7LPelVu5GAu1DlRRGAw0ocEx0ZTeGHNfrIAUXxY8CkDWy5i
LJczqZy/VO6vBgrF+clsdueqFNFwFcXuXLCKW0B+nWXmePOgc5JSM7gYpZh7Be7NQ3eEPXTI4i4e
krLZfKiAkvbfYbChOs3hcuBCmxA0+n4v3LPkqUi95hlfpobh4DwkYTjixaIxZlkLgzK19824l3n4
ke97AVEnxpaKWn2t6SQpzz5UvlmqtvO784ebFFajxQb9MTMT8yuqb4UcnviItKTpXeX2X7+Enicz
CIdmYkxB8JuvGDbcY9efTjSD4U6MG6KN+yZHLJhoBca7do37/8nqPy9+iDMh46d5D5qAbY5bkNOV
UM1HUuCIik//BXQO7NPAKaJxd0IHTfihZn3XaHUMD4Kr+4Z6hBvpORVmJDRhasomNxF/JIXMhzKS
tKJRdsh3QenCKljC6zoD+pmwj2Ub+sHB7Z61UL+giuVEtF9XGVZ5dxlf7Wepr+FIrxU1Mpp/dkqg
29+u0yWqS6Amec16uGgt2yqi6FDx4id8YXLntZD0gS1lr/ia3Ar5mNJCuHFGi9PQfivuWkYEWSHA
yB5XHJHO6VF7dfE2V3w3kz99LYreW37TMQ55RQGSnQcmINvvCDFMhw31AuNK+MSHU4IBAa2W8Fc0
PAuU6TgXNq6vcaNOd1DUzNU8NLihQdKigbANKWdeaB7D1UMhMrb1MFMKCtEkLFTB2xnuPane7Kah
w+OKyPD4OEbGDlcY8O83okYzdEX+iKUJNMZJoK7g2TtPeDRKTlBAiW1UCFjbHBEHDox9JdlivUy+
N4O2dsYMlVI8eCER8zyCatO3rOxNqY0yiZRkNsDO/0ra/CIlp2drpN5WGkYu2Ykp5YYn1iQMHyPt
/hFPZTNzxQRKmWq3ikqWh37QRBlSJjm7K34k/CASl8YkKv4tLb2lYn+D1J/5BUvUWQoUv4ALrWfR
nnJyVwB9hX6bD2PWNPm4V6G7hWuit8ifpcg2MR4I2M3mco6c3PyqIcwf1HaNgEK6krLWhIsd5k92
aKEgRgUo++PBVOa1mBu7mdOiYt4Mqt6ym8yewhy9Kow9TeHURMKiMQtpu9RKbUZqYpolUumMKJwN
r/azWny4WcOt13z+bl2aJFLJ5tU/kN2AlWl/ZjEyg2gOZLj/RDhXFNP6VhV4bxk+jS8t5fzi7GkS
qZ9pOUB0ob0sZsI/1WADUEic0DfRAuwZ9Lyz66pJ3mnZ5EOBrk0MZlR5S6pGzl9Dn4aO86XWQlb3
v71W/UGvYwwzkNLsTWo7lD9kyS4v3keuaDiflyx9/jrKwiJVRweRi8wG5HTO2VS50nAFSlzUo8hz
QfvDxecgzKo3Z+VZ2Qjiyfd/TVOg//cCTk2EvZJjFqzMHvX9ztxdm6wE6sDOrkWGsKKG/PTS4uvr
VFfLEyi99g6PXSa0RrC9SQRuaTRyWibQX+JS9myP0gYDW/bY4MidkG/yp4NU+TCnt2QawJUgir1n
IqYyotEcVAXejeHN8K6NJyvqT1DD54E0tzXd3hVlrFovbkZyg9iwgt6MUyj+AiEJCo5UsBDruHGg
xFJb+6jN74UuOJVutEcIFgLlWrr+gSeyTjXHKy1rSj0Y/WDI97odgy/fNWQDMCdXxLiPBf8AbWny
C1nP+DiqlhDdIq/qOq/oh9Xm5OFrAuYfVZ2H/lb7tUtaJDDenoRapRKmECSLh0CJ9oNQ+yhBjUi4
a3hSmJ3GV1/DAHaTTYCR8pwj5kN6aVfxvuQYOEqh8dOgg8Ule1bOiFYka3JGVe4Elhfig1rYtqBo
V0My2cwn11HWgPE62XUe8R36DhJWQkxR9rug7bDZ09sLyXUeZp2nsBoOVeYlHmxPCB6nYxoZ+oU6
+RsPHPaNNQh4lz09y4uJ2DZ/lJ1/MJJwBkds5Zd4P/OgNenuXhzXFjg8ewamOXXWISqgkTm/BsRW
9AXNsv46GSUY3oFfd7Vexg0eHjQRjwSfd0lqL+s9ZFFXq9myVAbjzz+3WgvF7C/+SX6Qe2qSv/u9
M07ZGsJsL8vbYy/0BcT7AdItB32jsIOUMXSgfdDHTdFdL6gNfUtp+cz33UfulB+PZO9u4ZMKAW7F
ax7PkFyuPID5uuFFlacKWvc3ODByGB2vK0qNwZ2mn5mCPUmAbJk5R/J9C9ID816tszEwUEsGQw/g
qbmVKFbXy2BEY9sGxXj/XZjRJ3nfjIHs7pmQCeWv8QZXplEv488vQE67ollLfQSY8uKTDL2VS38d
nHQv3gJ9XiMHXBfRLBALlu1n5/BEEGt6taIOAhlzD0u1cMCHeVqi6t+PT+Z4KrExIoXQKaDy9rD5
1SYyUzL9GyrUBlCps4Xl31KTX8R0FRZiuPawI0WJViWKcQtv9j7kyZsQFvwyC0e+cdMxMlGXmeK7
wcA1ObC6pS9lJWG89j8U9wT9CTwoKDRIusZx5c14wkX5JXM3eq9+vPgVblCK6jJr/B5vZLOYIftR
5gluZRKFQNjmqFCgv7iHH0q//Sl2vlWX1k2aLZV2SS5X3PDBxoxgqPI9Q9g+mYlXdOP/5u1Ig5Ma
H/tU1PyR7a6A6byo7339CWpUfpQZE9kJ0e50C5s2Qbcx9ayLwmTdkpsSIByzwcW9bXXCSsYkE5yV
zhbh+edJWmyhjZlECCNdHclbJXHzdnoEYarwQaTsJ8ZoiW5kLrxzdS4CCSvJ2ZPgF4z36KOSBI/7
DktYaVsa8H/qIE4mELQegoJxI030mwmvNBtq6baJgLAOUDxVn6LAX/OGWQDpU4HcisyqywCFxtM+
2oqXrC8zqiwYpSpCoaCqjsst2ing4IPJhavMOsW7fILcRZazPRB0eRnHq8wpLRj0uB100vWm/etb
cKibPSq6ErT7GIl7pRTxhVk8IEfnwDLH6BCKou66EWCKLye9wVnhZuiuykrjMTO4gzuVCtKq8cBD
gZPVHeSQ4hjM/jnPHJhDwSlcM3GB/6GXfm62M8nXWyDYFrYC0F8qfwT0nBMV/TZwqzmOs/7PpveN
aDGqg6xfDuP+vcUwn17p0kevUPoyWS6tHD/dDseXzBHTzGQxMYS29cLCEpd2uZ+2qKLW0GrD+AJp
5Eprqcg9KeHzkEHslo0i+to5iuDBU4CPdD79MP7QAKGyYpZf2DxC7oB9L8lNZAanV+J84Z2rq7n8
RD2kwB/2/71DfnurgfyywOXgfnQOXNpy2D6cTflXHipxJIsZe7OlmC0J7WvvEAbALHE0IX/6eD0J
rsLp+HYUnstpMLFdNOfLgpxgbQZHCvUvrD3xYq/IEkQq3B4cfnujdgn4n1jpMAquFQ7/e4hatNbq
48WVK63QfqVoJsnT06REguhoAu2/ZE8ppt2UolHubOFQMJV/WixDabkrntwep4ORO0ghABMGAUEV
G5mHW2ceXXIth6FvdBTapFxQbq8PVnHd/ad8JiuFS1HeNQ7apocmWP1Sajj7tqe8pqgASZx+jmt9
3Vo6fqLTAqFsCd7Tduy2egI/joD/Pt8fiTSX14VdFXFY2g5Y7N+K3LMRG6ba4PgIG1CykFV6hfVa
0aFS1+1yx0dxJYY97fvQuV8EzsLFzPD70f72ilm6R3rSBcPL8efKrLDbLW0wyVX/4SwKWVDK6zL0
fvp6Ca2RWEmdhqUQoNqjs7wSMns7eOXdGpID5qEA3l1s8ICUmriBlvnNlCEZoOzKaVIqvp6gREzZ
wzUojQhf32tAdaddu+6l3JXiM7AlvnB7dyZb2jo7yl2nGbJR8YATlVx23U0hextrzpOUCpOwRf5a
pqndD8SE0wVwGCG6dYgIc2RCjZjLCXmua9WTMktPIseLNwqzlUMmpuUDxVw6CGFhn/F32bJ8tXFj
UM3CrUizjaGpf/fW/zl0LKxGb6tVNXKz32B5LseAj75wLWdVWiidzXVqrVoXsWOljfW6DQ2HSeva
w4kMrFHDl0FYWqSo8jZaHxRxXS3ukby0SMjNHpsFnS+i2uwG2vOCGy99dyFlEpLoEDm8ZcJKReIS
S1ThpX5bLqV+wGTK6JQTLqRcnE/TdWp/tVDeWBM1eet/XOwDiESDxjmbyrxOWTttTOd7uDeLJsQi
3Cgg5bBjDV5ptSAmRE/pjNxwYWeVIWsnIPSFMg6m2I2as0W3X4d1fhaOwN3rcXZg3dVikHaddM2Z
Mhr++yxvFS4H6eDdwT9Thx1e7SVnVWvaxXgqYZDrx6DPNtS2gG1c2P7tQGfikwvUVl0nd0tTAey+
WOGwsi7bNBuDkbc6z75pyzalSkjdD0BK56VfDjOHwLP8ChEivxlj+Kz5+YeUh26skM+dEJlblSeZ
QXaiKG9+F5Fy2r+rDEvSRlOGFQ/NTw+3Ks0S38znx2RgjdAkDD/PPzdlCcB8nD8TuOvGflhb8rpP
9SwGRZVMc4cwo85MAB89cW9cI6TxiVHq91gqHA8D8a/8UjXFDgqJQA2IWoonz5vCTTQMWWaE5oZO
iHvct6EdVumEm+n5i4NLGEm1TB2ntqUpdRqwwv6ZJkEbE1DVP4k0m+b8L68HtaRCrtsupIYBd1Wn
/cNbZvi6Uz8yhB0PRE5s03vOg8YLCRPPrvrFeXMjTptTYnutknNNSzzY7qG7UgqJyH/puRVNyFD9
xqbBptzF8AZX74KRf89CBTCmj37pgu9RatukZvaCcwL+bkkccV8GE0aTzoEl/tS7zEPuHCk7hto/
uLhZOozq0ncEegXxqpzOS9hdYTPJPVbmVDzsEgUbh4PeMeRd0F02SYX42TcX9eJAnxEEhwonugtF
xQ6ohz30Y6WGqTo2h47xoypvn5LE334FHZ132AMD/vlRBmbUkyGeysyp1eL1Q0g9YJEHs+52m0n4
hJFr71hKa3FMSkFYa5/UKLE0gIaetOQwVb+DoWekQX5FP5mB2vOW9AfIu/b4jsUXF2hEdTPahfk7
W+bKeIUNSb8H0HdrGnh3dDEAA9gms5xErhjjeL0eZFflG2BmaCK+pQw9nE1rQfESOVpQWzQ0Om+b
O3Mg0looh4AnRk2X2n3es2PKLzm47HqMmQR0x1frq50LCViogdkT/5FupzQqbuAJX7UW/9lTMyPJ
hq5YGXatpGrBy9YSbbxfhZIW46d6wH+ZP9xXLTjvvTl+ggNGUYg08bhSku5fDFapcwX0JkKnxoEZ
DsYW1HteCewnzZSoXm6pDBONi8xS7cecStSIm4xoKeucmiJkkKkmqfPMoV4XPQICvYr+/FU/i49F
/pddpkeEbhHoKKECT259mJLqcwh8S8gNBUiGJdqUCHijJFe88Lm030JH075qYo95wsXz1XlyC5jm
Tix7GoVR1wVbEulRPSWFg9F1Iu8+5pb0qODRmyhEdLTAyOELFH/CUXzRge9hg6nXrwJLHuAms3I3
hxz5a80T8KA5YWTE651RrGwE8L42eOnf8wmSOgJbVtwKB1tREPQUB2D+wZR/UqetDFOZJtXcuh9T
/oKbT+aMgXMBiAv2SMBXXulMQfGS2OenbJukwNsDPwCSciecbtmXmoCTV/LQsgB4TNwHpigsD1bM
MPJULHJsjX8aosqYL/YMR2RjirwjjrRMCEyZODbQ8MYqLPVGlzWXEqNfAooJwZ+ec9/Hsh52dY6q
JrLeTMy7p1E++I9ts0z3Ld6BpmAKOMhmpEhWdvZgwGecT8YBhp021ZNjCJ40j3ByT+2igr6jM3nE
PPJ+jBKhvhfZ+gRl54Uxv806aZYm7jDXBJ8QJLLXGh2G8BJyKq64tMGxprleBDXYbXDytLaMQX+c
RooGy5ZO2T/7ELIPe2PfoxSjxfFR/KoWQEPPjvigD9+H3HyCQ1OJQWpo74DkHxVZjTpde96OTxYc
6mIchZiG7zMMpykJ7qRlbxHUGEa/jIXYSr2M/w3nwjza//qHWJMQAEsi5Yn0x3zH9JsFDqD1Xu1v
uldihu8VsyhhvAHGV8d+MXunzVhmBSyPEU5BsaSpU/Bzov4UJkb61Zm3X/ox/38THgZS/1j/SXYY
Wg66wFRtXNflIrFcoxhM1Bz8aqpMveTFh4FpOjBVR7maiRS4JfyqKsas3gGAPPKdl1dw3T2bLJyQ
OqQruP/NpY0YlS3JmnBExLHMLqvg4MzTViDNkyxLV/V7uNo9ujaRiAXeGOPLhJmxrOYj55ABMxqz
a8aJIRZL9T3HxxGPRaQYx3F24Mf+NLe29C07UVzArfbjA5PzCoKq0CegRyZqJeUufRdWncIQrZ4h
xy+BOg4hAN9QYWZ5yWbX0E/f2V4c3gJn+QsxhAoYYbNS0wB2ndlQXG6v8J4C8/TKNFDKAvRmKEh3
W9Y/47QIAudDOBqb/TGQLd8QI6hdoLcvwdbcaZ1cl+xOjwFrZC5pQ+JTEwP3Jp/ro86TrIJ+cbeC
8XhcVl6lHhQ5hDxH4ffClKuRaBxtAgpfHEFceSt/GOptfN/EW6jr8hesYf8jYspbauDLex5X8X1a
ggx0lwaEp7nMcwjfZKsQyV3xh0ZCw0tkd17emSnhV8UuR7MJjqUvRC7+lPOu/gXsqDxXhUvLmIrv
xgq0psiN8kAEiI/K57RcMI0Ic2K8GF8sCoKENa0OHla/GiyZEccHyAMJgpmckW32mPjN6G2cGdJH
0D8Day54jp3+4G00VRQeYr0gjIzt1g8Yz+iyOfYYkt2dBCv5q6qknFvqKgWWCBWXp/CuLfuHiLhi
NEfB6WCHe50YWMHdjuV2GwHsK9mZ8PECwV5xxYNxtRjxHoHwHk2WLUtrVY3qgwQnh6VVz5N6PwbW
rQ2YGgEi5bpLH9lrnmadWcu+9DQAqYxrPh9cX7uAI53+Upi2/582bEpeP8hh2GazYruK1VXoGm8U
Q7A6MXzVemSh+0KqHDnN4ckoaixU5Y/3dysHkIl7GKuTh+hnwXxmuhTnuj4jw+SG+5RnOS6ym6ol
xQ9nQQY82ED7Zayv/FMDMFk0W0BkeuGfn9++JjQ9K2pOr3atuIMXXewVn+UCYCG4uD+o2Ua6qKtS
bpsUDjRZnP4TQXxID+6ZnRRd/g+2hTZyGjWIahsddhWfvInK8HXPeoVMzUynHAxiA+ZtHDdaz2OB
nkIXtFG0J6j2mdegLVUruClmtd+IdKdsMPP0KecFs7ZCvNFnyRFT0xHwW/OhYE1zjKEvagAbTJwx
/lzaSYi4golADK4Cdh0T6YT7q0qe8biv5BMma0tJO2jd0knfi3e1IacR650zVvlbezVuwIxbyI/A
8QfQEcEiAQsg7anivWWRA5fDs6shbWdvM5/+bAJ+HmsDAHmxkgs8oguYCTzbq4NobqAMlXk3xkX9
Kfb+tGNz3muDjvD3jpBjwA+Gg7fFWr1j+ty7bQW5JIuaOGRY0eW011f5Civj//0UtfRfrG1SZSSg
sz4SWk491nL5xvQ/aroIVCRFRYeCo+X5kwWC6Vj48/dEm2/mAsMWg0UaTWCBWgcdNLVmukjIC9Lc
9nSfoESTPYVIGqiIIFLduGDx+Mr6vn8RWXmMgb8QgXTsACrH5kflr9s3lI9xgokC8+0E4g17vkN/
x23n4spLDNeGIO5GXHH97bMW7sISBOiwoxAWnSLYq0vEYrJpzAISh5Qdt40eUpPyyNhdx9xufO45
brDWI0MtXVmaUwxQDr1StaGak8Pqepg3njwvu1g/i+vFnc8azvvsEt206vP1Gj8QG+pcCagmEZhK
bn2J+JcA1aQRF9+H0S69J7n772+01Z/QJuqGwuF3BpnwZzpOFDTr1PHnZDOZ26ht8/HyV95ANvr9
gRv8SUPV6P7HVGjIoFUW/VbfiFarxZqYuoxbLvOyIE5DHq6UIgXbCeuG9YrSwCLJuuNrxvADKvm3
a/y2fRWKQBDCrReWkjBS9tw1TMwaDSyZtjj/6mGYRG3yEHxDfqWIDJmxjBHFCSftOCpvy0qxY8iG
TAvdx7wzBhq/kzPEn2fkm2hpEtEjDKYhVeHl3uddm1wDZQu+igxl+8tRzOnAfAO5uCeQZD53cXlL
/zznYfyqTgyr97OgJEUCr2sv/vwtNrmjVF6jbO0bzBd0l432M815XCaiqlUkakgL5Xu6cratVwgy
A6ewjw+mCST2Jta9X3VtAGXex8ydrypJcESnT6Sc09cyTSvtvyiSamWbY1xQ6PGLxyNID8/2HbqD
1KFvJzPjI1+aSruyuyuSxhghuxR7MSa2OemtnydORhVg9zYWPSCILcaa+rAsJLyYT2PJPB3hb1Kc
69bV4V+45W752oeN5XSrBs3PPsfsXuMcw16t91NeyUBcrbYxD327o5SiywAhdtEII+d6cphKDj/z
7M9mT9O82LRWLCiuLtLH0udotnjwOyuaIezwFRVRbQrSAt7W+BEm+WA+UYxJSVGFIom3Ah0N8Osv
X1cu/4chIR1ChI+Zbga+h4YfOV7TI38YQWeBEh1fl+3uNXMs6UpWoMxn5daKdVBokq0Udk+FqOPb
Tzm+dXi8+dJIOWCWBvbRQVHGbPHuqmV5LjVB4N+y8nAOlJlBAbMpGAmbt4JUKhVtsU/Js8nF50aq
fCCe/jubBRbLpd6FZ7dU1+FwQAVewMfOxiWFwZWUqJPtS/mjmEr+02MTU6asJG61b5R6v1xdgFU5
Xrf6bjn4yEO9h/JN+N+CCU0cETqfezrP/YhlXKrUiGtL7XYgk4mpEhapt7ufZv8GkvXe/8K335DF
V1tD8iCCGIcQbVq6dEtpMozPUyHHYY+8jsyPPDBkbMuqOUDJykmdtaLXnt0jGoexpNl/7urApgbE
T5zo0rvj1uulheHdujl2n4xX7QCuU7rXS3mkZ4TpvyCZN5QVU/HN62kNlZSOmiclcwkDD4IcMO7E
T+YPAbEMzAPdBAlgBUtI+ZsSisePY49P5bubxtJL/mCRxInYp2Ea+HKZZwSMV0ZUusrgsalFIX6T
L4HFvE7O4BvqBP+qBxyanvDQzwfFSTP/nZkrzNhaU8GlirufS4Xp3RcNI9T0EnugXGoH7ND0V5La
Svd5GAGP0wYp0s7+zMNVhA4eZ06NukpKXwoL5KxhYV0RvNEhh7Azoi3Nt5Bq3R763ZXaQTrCtz9l
XI7dhCukVxrJZV22OTcr7GjCtxVwBtKlrPuQ4ZSQmgchqR2aQIeZNYeKzMH7hFl/KsTzKcREo2M2
NF+YGpRtKl2ZKyFqmFNB0MJZRFK/kozn8uOtFMbwSISF/JAzze3Xtnkfi/9IWlOen8lEF3BlwF78
1YU0lfqcr4JpnsUDwuB2A1z7Q6pms7VtrjcrIPss2eT6YnVfXCr30f7aN4Qm7ect5VdsPXde3pZ4
XkkAyjUE0JQOYPOB9GEg6YaXVt6R+JGdzNJeHlLHNeCCTOsBdBZJc3r1CyCI94aYt0GMzu9cBGX9
fQEAJ4+d9Vwi7WeajqbBqOxdON1QAzcw8qI3ejIkR/CiIzOD2V8Kq8q7hPg1MyK1MyYriKp6i6EU
JeAE7OF+RvG3h7155cy1Dcp9uuFmpca6PDgeijVMNrtJ1wwZp9gEpNWaqhTWgO5RVqd1wvZSOW+o
ATeG4vKxaNnZH25TxmFXx6Q5GFHOMdaqly0oguEynHnQP+mWyFgIbbydLZSvuMqtQnBIJ3Qo1krM
MYaf6NUcSu4+u+ki5LbfdkE+SkgBA8BfSFTffdMXqhyZqH7r7JsMfEtZlPBcWkxAROuOFo19McGo
vDjNVBFiH3aQTxBu9/q/iLZVgzFqm8zwmvwkPdbfrT0Cv1P/K5GTPOm2Ksrs1LHb/5nHnsixzpD9
K5SfVRY6mCzwiwG1MKlmKBuyVByZN2/mfBeguBHPWZ9YyAFqJk8XpUrMUtXj8v4Ik+WOeY1mG52c
W2max8K/AWP4nHeC16C4WcxLeFnx/PKRXwXNzcZheMZByaWfThgaTwegvMUdAPNrW8O66UlEAy8H
cdLgeWcdG0BgtqjWkkAbft4/pzhSrCapU/imLHBiiWRQVUJZ76CuuFzK4M8P6tXOleZWEUnlxGB3
NG1JKObTE/kmz+k7fTVoTnxML5thGjwadEp/18ffBO3rQ495xONZGh1Fpi5TusdpCnX9cCRc132W
UzrBnCCbhv6I3tNaXtSEo36XSxpHz/654uO46x1e6l3xFt9vftrKxK6El4bHZpKmypmDbcN33AW1
9yMS8iWGy9f4kkU8UVRQIgdLutYiJxXiWsXBi27LZyEZ2JKvbd/ADp8fQKf7863fNNHDGWyPLXDv
TRbYDJA5qWI30ZAxoGmWNPaNSzaEg/yO1M6AjjlLS/WWTORCpgy7ugBuNJPxMZzgE2lTfopVCHJK
HN5mJ3EUL6CgL3+QGSry5E/YHAzGs4YuUxiqRF6lQ3D9GB5C08+RQlCkQfo0HjYcRinXNo9nnaXq
NI7I+WawtrMrvBYnqA1be3iUiBcimtAgINU245sjzYjHanizmDCONRVR8bmZ7/8AG/MVGMMl6/zu
MhytII17WgwmgJT8fstLRCOrWm+4rfwogVSFwcFLVz3UZFUMF73SvabqmsDLMC0PtRMhm1XKZYUh
pFuSW1bXuxXOL50TCIYeppLKCG4wr1IFsd5BzqQoagVBg5tJwgFo3SiWfXiU57LwpZjyfc/1lXi2
B/d+TDFBnMn3brjjf67XYwi5VD0Hv/DR3t1UTwULHqtVov/KniUYNzK4Lss5MibvAkoTp+S5qQu1
tm3BLDlylJs4XAzTxwnoOHcYWEsxF0nm6efLPoHgK8DrohO/w4JdJ4NdNSkbaA1nuMAbwlGOu3OA
BeaBGCwBdKIr96F5Q6KjVHKOqIKM/epxRXpRL4U9YnZeYSZjSg0GCl5xSEZp7+r+j5v8HfrWPMo/
ZL1y0dNUXrJsk0T0vWcMWc/kaqRuOt3ahcMoAMtgjWqVVG2Eo6px4hMOfoB3E2eAQhgSlUwIRcqO
yzLI/0lV81NTL+ReqdN1JtLN0+sXojRzuwJASqf4nip8jvyo0rvqLT+SjPU85GzdI5DA4LvgVukV
jdMQqp6a17dEAVthoWoqSdHtF4WFJwW7c/CuU7SI27rTcdQnsqrb8/3EpratzI0Ivhp+/fST6T7O
4awxtTd/bQwhDdPmqQYMi6xntVeiRED9DlKHTAu6hPP+FUVZFrFyX99WCl2L7sKZW2LE1JJyoyN6
ygpgk6FHX5Iulhh+oZxAkbHVJrZfc6pBjVjnH46qfB7K2CCz8dPSvvYy2Q78L7A2N/hbaq/3rCqV
QKEWb1hTocYmDaS3F/Prm/C2Aj8Lrx7U4Qp5pPF3lcK0/4Jg4OYRTMVDF5gQkyDQZ49cRfi9JVpy
m72Y+Ks6GyJuHx8jT4C1MI80Y8VctrXb+jDWtfN1XTDZQR7O/shX5uTjHdlQvGZMV5YZYmZmaO0K
KTbrUVZA30VLVPx6JsBclZ1PT18vsJjqSWyd3ye4N/n5aKbs4/GDdaD73avaDUKaKqAHzgITrJKf
fp9sn+4my3G4aAK47RDHu/EQa5OVruseYYixiZdqOzRMEkzAcHT9goktUsyp77poCJHQrG9QxBUs
lSYjwEyIp9C/g06dECGAfToFwJizHmBk/fCOCcEC2Z6hGDMazwPfop9ZJnrcTeys7gLLvDjMJed2
cjwDk18rXtH0wX5O6+3hQkKC/xcIJsDJIZWoWNK6xktYklsg3v9WiT6wZOkyxpa/zLwkpb9oxJqd
8SrpnXkwQCkV/gWMG3KNEqT8XOcOD9Jm6AVp0ZoAAPy55qh8csJo0uStUCFAPcq7fJmbXDxIyxmi
QYRsTFky+bgdV66bljWiGMDzo3uLh8k2ZYlldBUM+uupFjtrk6mBT2rB/b2Z6wcLhO5D3jOF7xsK
G/EZLXXrkQX9DQMDTGRBCCNrV5BagnbIFM6IvrVPRS/7aOwujOgti41436gfzC0gZ7orlxajVf0d
2duhPYB+/10DsXDdrNxJLVa+mRMbNuHhjqZJGXzWQewt2f4Z9Zv/mx/VZ/DtmVqxb+KO/uoCa0au
UYwEmqI1mKeoiLEjvKibcn0LIZqMGK5lNE8Y/n4dhe0XPjlRA9QSWxbU1pAh3P22fPRs9Oi4Bl2c
7fwdrm1YeDE6Pzne79rGt1SZl19g1WKMq3dQ2izy9t8eFPJoMVfECuRoBxo6FgwG+abLC0TcJnl0
Hq1Sy9USiqjMRECprqkzloVFCliMOSt+PlQmSFKT8BgnogrZtCyX/1uEri5exvsGmzbkW/twJJSh
l+D9G39hOWw/gFVBWVjVILoVsCz5kJDyiZYh5swOXu9Yqr+lBt6X4GKxiTgXlVrnO0St5UC78xar
JMRau355ZCzR//DhA5vuJcjJLDGN0tfKb0WS+NCRuA5zA2qR2h/NAP2h9EEOaVNHFGsGZiB7CPp3
nGjItY2GPqG4lWFEEDoM6P3JHhE8Ge+L7/IIzYoZRyzxyR5p3MvozBW9QkTterY5I9oFIcZnbH38
yS0GV7iavu4S5pgJNZENgdwmP3zdWVAe61lLxb6nKlR2/fB2vqaKWkyHj7K0s8C+P31RgWdd6SYR
axMbdN1WQhEczj/fUUOTqw1Zo4KLtt/yEitpFKSDxTS5/1SLIk4/ER8uO1sghA3JcwUnj3sPMq8E
u2ualGa7rW5vmE9bFagazjWeZYg+g0v5BANSWZjvDIf6xc463aloqDLxV3G2aTRT9lTmBRJKCuoQ
5Lknpm3dei2A1mgQy4rxf1jwK2uNCpueF+2k8HGRPIbErwDQnxa6evAY+c7XxpUUkZ9Itwl7ld2/
4nonZwGNkVZYtO2THM42epJtsbuM4ockvteL4fJk8PRfR5/aRhiBMgtjlwlelFDDpnCgI/dDOFL+
M4rhtVeA/e1UGlVw9zvD7UkIEJ0J/jRoQ8UaiDSkTSd3K0puABXwn8e2A1zelXXp8XarX9qY7tzB
bZcef0iV62QJr0FGYIeRahEO7Dk+5bJ9IeQPtOdYc46QZbEJxBUf7jqC4FU68TZ5vq+vUZ0Bl6/p
cc0nQu+rA64wF3wLB7BAoNGqz2rgXiW4y5f9x+jSFvw6ccG2OVl8//mU7CyYyOZmU+p5I2x/ou7a
BKnRQt3ThlTS1sFqILwrhuvW5iFkNcRnWoeimnvSyQMCgLw89DR6gjGJ7MS/ajoixGnPdjJmFEBX
UM8EEHG1p/+IeEuQ5ll6Mo+TWeQFQ8C4Goj7sB8JBEesS2cpioz79Ot9STnLiILdaGEj2T9uH/4d
jus5s6P9b8K8/bq3c94J8HBp2ReqhV7pJ+pZ5RdIWv1oKfPKCKgvR7LUH5zthsKkzySnDpW8Y41y
QT+bX+/aJ2RoeQCfze8h4DEA7+WLychcq5xv9fRhbxsSVLeKlHzBNLwuUqnOhQuzbSbwGDyANffd
PhpXdAWPsdxVjYPaUhgPCmDBDCnVVCr386CHqYhYstCe/CUKZa9HXISO7vKUmGLkimQQIa6DuDGA
Nw+zy7mNwaVjpdH60oAy7569FIQQ6nfL7XuNtAkfwxXuRFBk2r28LxibqIMYAxsAMKenehJ3ageT
kto5KnM2STwoy4j9DFYWmSoBioyXbXxDwBIMGEeqDWCHo7ChPTaOVhbS2IHLX4dznNk7xrAOmat2
YRJP8q4fJ733zskvKDYShNXbMElWVLkeHQA/5lpoCKAyob7P5lVCTBQ1meYcShPOhdF4gH8Trf6w
YWjoDuHrTKLHEWUb/eGyIeCthMDZKpngIaS0p12zWWcxT2ioEM1NDVlFVhCD1+vyl30a9s+tPsfj
5VDEzNXOoiGIv2IYFAu7OU/mClaVML35Sx4qHSBjOgzxx9OsCCYJCvmgZByqd9NhTwVhqRwabiqm
bP1Zxl1LgLeiBv/DC8XkIq9AA6qb3Kvxh0nEHV6eUO2kStodRSgssbBa5SO7HTGzPwQyZnKA1MuK
HQXxEfN3O4bnFlpBS1RFSWPhVjbYYmA3WFDEtESQJ7lbHvubtb66Abd8JvMN8VKgcNduGE/KegEn
zMpjx3sbi/aCkRcTyAPS9clRwrGuG5plUGK/KWohv9ZXp4sT2gOqRiCef8vDqYIMS9HWb+Q8igYm
aUYHwu32KyWzMdCrSdoroBvTOuex/zGlPU/QOlKs6ndTokt1sOfpf9VrFkEuaD1W06d9EOs7nYGy
1suQjYchXMnu/Du/jPvLZiXCaD7qsTR/FeKylOODWpKGg+gOWGZHzTHeD1T9nxvvsuBmJyqYI96f
QchXNWJgAxZ6nGWguURuhkhpm1v4Kwl4a4J2zWNUP86q9nLTh2b/i0yfm/xf/Wckrg4JWmDNSYA2
wlL1Oq5KJGVY9ylFDrK5mrqGrAO0akI/TgJY90IJqQnN9EEirweuEMC8fnMso4zzcl0tXJFS5lRN
fWapobMRMqT5Z8Q5Fc1afoO/yiQUhP2DFYJkFQFyGw9ObFZlkkQoLSDeESuQMqayFqcvQSv0oy/k
lQJLHbHlUhCskiVpp/9qJLp1XelgZv5ZRSQxFTmGETI4kAv4tYxj4+hvtbTO8AOgJ/mYgYY2+wHd
Y6WAosntsHTS1hVCQvoSFonaeeKkSTqMJrbcna7eVJ5S7UaJo8U2DgxwD4v3Wxp7HuNbXK7rAP9o
u01jXUmid1iLkjqeKc82z2coZxL6UCHzcCHfnflFJLvCRFZXdZtUuw4GadNllCBXdcL5SCIFdKpe
KsIPcgti1U+DbujWNd9Eo8tWnK7GUJE6Pt7Kghp4fUZhHb0pbYg+4f0RB1AtyIHFHWhm+8ym+2U7
RMpmHZQTLPJh4fWBlgzidxmK/FQoF9joF9591dogFlK1qEkNGMEzejiO4IK8Xpvhc2hKgfU64rfc
mCGnw/VqoZG2LiJr0SVUzYCH/gY049P3oQ3nQAW/GsdNt3avo2k62mEoJ+X1GPe9oAACtzFKBkUx
taG0pab8UIeOJpwJILsR3KjPS4YoCYVuDwaV6n8K+dKy2XyKo8iyGZxP9hBp+5itEFSmHDB5E8eN
oWzOhzqe6QvhEsOL2O1oHvBADjYIx4lwUjwYFmsPK6lmXTif6I737cSvNHoCWJ3BKj2CswjXyZq1
HFQj+tsxmJBqUzSUv4wGsJ3dqlbXeupJIiL9RKHSrTcw0nsESegi0bTytQcexCtC/JIyOihS/aIk
Drs78T2DK4fd6f6BA+pPINFmAxX2ilxrbPbDWuT7G7GvKxjF9hjQV0jdc0FoPVx78YPN7As5Cq8v
ezafcHhZVGUYdAWlvN5sod7DCgGbuiLz8xDhSPSLgZmcVT3R7llQaJ9IPdyTqes/j4wW8hyORYk3
5efW7QMCTKbj6xtiOER9//1gXmDj6gmFEzSzuFLtRfR19lZuC6LfV/KiPGd06IFmKbT06GLZSZZv
sQlXMOoeTMkAgu9OUOr4O78HX0V3USlU8+8/JLjnz6unbR9aodfSRILV2v7VSkrGipiQGY2BSn9L
Duo6NQyOaPZEg1gxomM5d9gWXzuUtyJSM+5SggnJA4pUZl0irplPsLGMR0s8ioN48iSfIG/kaQi0
NaCE/SdWGhprpkBDpNoZklsoTb3sPkhAmys0o5y2h0pLypbfmw782TjaYSmLlDrjFMCpHcKAApZp
ymFAvcSU8qUJsw4x8d1+aDZp3XOK6uI8D06VzoALxkYZDJlcqOEx71qHLulRE3pXaQ715yAFFx+h
Vkb7kGKrhmQ0Tcbss8iKsQSevUtxpjZeZ5XvboS4GpzSO2/LTPKdoNiejSqx2XqwFF0mHAoYEs2b
LMk+L6vlrXhkyaQ2+aALfwZpXKTW4HUzpkExq/HAqvpqA5Wc1IHuB59s1bVdF3H/3UVq3jxoxxOs
Kz2AgaAXZo4F1lvkMq9blVODTG1yWjK+AClEK1kbJzMegwQkqV8NweetAy4sda5dVmsDa+gUUuX0
xcwdxAJX/NYyhVPQRyYLJH7o2mDxzI4nm6uMtDx7YSdrKROIRZvYOew8QZlKsuP3wZKUVhbtkSR6
SVvaHmbiOzqU99ZwKvAnkwypJtP5WWk17bZonfhczNxe8cawbJmoW0H+IxM6prXpVO3pGzm3WR4f
rqpQW2whmPmvqOvy70R9MucfnLuDiiKQ8rdWhzFhyLIqxui9LFMICwvCd9mCvDNiL2otJg/hLqmL
j8IRCHQjNocg01BvJYd6wx5GMz38RsR5gae79lFk23226yX//ZqvRa/fl22NAl/SNMt6m1mR4/o6
LsQTpEzuLdVgaaWzhgTUS/weR4Mw0mm3NV5ckSzxIR08h5xR7RXIffY8zLlMIHM6JzoBXn1bhnWn
XSUw/AZVuZe8ExHkjfRI7d62hsn76+X7+k+PW2qzIL+/RhePd1ymLqQauUQHYzNGMb9Mr6681HxW
oSQ0nL8qLuOOXM0msJrVt2Zk6AddFPSCg/LCbMIx+qdCBlzpXNxKtAC6yq5WvV5MKv+bOCYfhhIk
tuEtCYi/ApFF8/xxX+uSigAKJbyYIfUEytbm86+DCf6YC2pDsdsUxmbotNOUMwPtRFh+W+a1tAMs
8DuLnsz6o3r7XlsP2703sDFzbvOrrZzEeta2U+/itYmCFeTaGee2tOtvW9IV99LH3mSPQMj/GTzR
kB2cx1a31EZBMJZe6wUyj5H+KChDBVJMBhCWFNFQ20YhczkTNwJQ4/RKEpD2+1alNqR6X5G6fCV8
SBQF7eXaQF1Ve4HSfnx7GSehgNjIgnLudWdaatvDeGSmM2bbX7A0hsYSBavid6QRU2mxDghyxIUc
HZVlw4IyxT0MNH4SaoC1VDXgNJIQml2YgTLw4Y2HmKOuD+UB3Kruvn/fD6su4ZExfC+1FPh/2JwG
tfNyo441ntSP55doOkPsiGqmlPYLKkvDhKapm/o4phUKMmhe59RbOP9goiwj43BdwRkXY93RZL8n
0daotmR3CSE/QT1oJSFTU8/bhaLDf+DjDhyHRQ6sLBEf1z/PN6pCII7ofDB38M8RxLeDZHtgmQ6G
QtKWc1T61QRRVQJ1HMDPaJfQU6uxDoM7uUiEolklUE12uM2gmo7nbDMXI/NUTEhA/3vTqgVAnAgx
MIiYwQ/MZudHlYvP/qPD87dFTjiLo2MXWwHt5lWgAejMkoIKBTwpJTe6uhghKE+5eZRR4TMuC4wH
GuT6s2rfJwRs0WHsXS/1axqUGYOWWEfmJGtGETfLPl7IgN4A4IfXPA6/zVSXGbF/VxI6TfyV28WZ
gsC8caNlR3EnsXhxBcTLR09hEs4Ek3BiSYZXDkbRVhMVWG+mPusSL4ILt8KBU0V9b5cNZv/XP+QS
8b7bUU/uH70Wbr+UWA0mGiJLgty6pDnPVJ2mnqiw6t+n58+VPpE6/Yx9/uZnzJ7tncDQwLiuQewL
Ct9cuKqWapfbBchgazJVv8W8XAEZxpxOGOaDre3F9zrOOH/XOgvKA+IjvoVDs65H3JAIe0/5ro7l
33je7PSsJt6th3G7CU+NvTrqBBa7S1MJDqdZZk/IuGjoFesiVx+StU+ysyIo/IISLeaFnOOT04w/
WsZtKMDw7m5CGOrUbd0Cl3ABXTWjeMpskmP4bQqD63P67+uvtsQMz4QVJ6iM64xTz5Metq47TOuo
jFnN3U8f2Y0FwsxysbFr1i4WBchpQqOCrwBVjoXaODwdxshtvUjF+V/uJNzx8IwpqcqygjnkEbC7
fXFDXGZlluTGwbytFRdYxLj0GKUjHw52K62wQ0xiiizUP7hFD+9+Srx6n4N3Qdz6vHO21I7sME9B
MEkSDW1Hoq+MENmRBJvFCr6vltNjJw9rdbErBjVxTbCZMvgo9r5gKttbezu7l5+kMxem0YUXMXPT
ekKKeLkg6rcCi2EwN4Bo7ND51Hik4JPK6j9SU9zIzLygSip1SRf/xIAfx4lBK25CzyRN58xm+LQ5
zIhHilQsJB1xf3vn+JDZXA6df6JMPtOhoZt6jrZ/6mNNnJb7SsDcS3JhMjlKI8j/9XdT46oLNpbx
CGAsjKbq3YV0qQ3Tfc831AN0FY/hiq4DiXykz8UQWYDzp6AHJ5D13ue+y9vwpKM1ERNPJ5fOp+Bs
ZQAQGiZOIvXyruQ1+Ydh4JCO1LNRUtVm550RGzEN/m7pQ27OcvMO4ZT1pBBPOp4VT+zfaKW/vNXA
xdbGtZCS1ytjDxbUZ77EqfQ6fSKzNFkWMP5F0oPxOipzK6FbkPdduQtAwNaNWVbIHYdIlWmomJFF
7DPEY1pkdXwzN1ve8PMTVCbNCKuNsMdv08zWdFMTV7a61Fwp30goA5Kmz5uqjWYxM08Vsnwv1Kt8
81bMqa6I52LRJypeffHKyw2Z/hhYuXks5kaBaf6hvBhEtX4xt0EN+BGzJUEpaUhm9dbylsOh5Z8L
O/myTdgqtSQ6O0ti+L3E4h1DurDWom4S1Q9q5VjcyktUNeNJEh2Rk70OJ1WHoZIisyvSy5JRSZyR
TOgeLapc8oLrvtLCeESkq+syw+RqR90oCVPltSBv2SkftDGx0zDpv5wrsHOmB8LZQznDEV9C3E3g
9MV7NS9Veuq0CwC/yvueutCXB5XSDqQ81abaYeGxbJJ26RucZ7z9g7454O/00Ktmgf0pegGZsK25
7ylA5y7yRrQlEFSAXQHcX0oInHafyo2yfRsNrGrO8D6UfMmUnXxZHgrorfEdDnDqf0x4mYzW1HWv
1+ZwGE6nEm81HcuHAhlGccUt0Lx2v7mVWPiRxFQWmUMRin6St4j/VlQp87gGReUkezGto+94ti+v
pRyfnj/fq/YqfkT1PbPQ1ySSahX4dF2z41eUVFynPWJOQrmR2Wf0oiYCRx2eyqdISqFacRSw6xgX
DUg1GF7SCdyw5dkSwKRGWienwIu+tItMxpwwC+Pq6A8ASKSjBD0uqpWkjaL6FcXWa/skj0SQvrTA
cRbvsPadt3mO1RNOngCbIig9vBcLmAvWq4+3koXNTfguj6esbU33HIviGxE3fCrVnO5URXXbuAdS
0ho9+lGHvLbKqOU2TcAMDDqma58h+Krm4Vjjy/1aqkvww685zAg+upgoTad7ywcB5vR4MwuPqARB
FMMJQZi3ZUYlo31EOurY7w0OcY8zQDJGs04VqwqsIhabUsUh9vfDuW7NebOWLhf2jC+dxPBTp07f
HeAlQRx7wRPmC5eu8zgR4FXTjGKpl+C9vdcDkbXRwjH3ynqSWQcN4KYIJa4sPMR/9ZA+k2kix5OV
ApB/6Y87FQWCw6UYfWt3kw2Uez0WDylzrssyhCBuSYW983U66W6ROAcKAs7V2p8UCO3aLSb6CsxM
OGNOKa3hsFFAgk184Tx76IWYqrE3gyTp0WyjinxIxt6hU49ji4h11xY5+9KcvFaB8+SwQnYcQYz6
OLiLVyRvbecwYBJZc2aoGrq0Lix9sw0QdLJGp+TlDqyEWh4cOtOQz14KjrOti4RNTMgymOmVaUFg
/4DSrwR3qV9JnBaOS+T7BKnsiOhVmSlVzzfpCWL3wYe20iKc1wl97KlYtmnhhFwjKGEgFqN/9G1X
Ja7r//67v9kjFPZ4IZDVaaz8vhV1NArwHRzH1+0Cq5HwTgAz/h5N6LyBB/14uc6Zz2+OjB1t52kx
DsVOJBunjugseXZeeie59JLJSVnUeUvxDl7YlWpN0i4DT8kALu5A/zm2viXXR2sw9G0oiBaLVS7x
tAe1pUJ3WSs3C+nuzEckSQpGSas1Qj6wTUWWtQX8cqdsq+eQH9eLY5pd0z7os9qDuBd5QPkQeCEH
36P+xzBL50BSq2nO0are78tjoL6P46Xc7U8rNriAEcBBTWubc/Q6/5Sq0EPGa70Fwp1iIyv9WeaG
145zThECNLHs/itqWxd8A17D1qlCm5uE5DiVgJIWljsrOzB56QKPZkfseiRyXNm9QT/HAbLuO0Fr
9KYlffvx3gzqroj/CMXpmzubpWlTFlROFhfLLJI2Uvy6yPDQhiQuQO3xuXA/DsPd++D9HQayJImm
sCc2SOuFSELDIAo3ku4AtUv0nAGv5o+MWLSsm6EE7mmJdHzjg7xrbeH/ti7mMXDBdhWHQrbvHnmr
MmXQfcqVgz5BjWsUwmy6nN2v3ohFxlOkxEqsSsQvqJp7jCzGlc3fnSUJpvNc8feJjlAXuB7qC8e5
m0NuymG1inOYHjhL6bFLBFc0HM0IR8QfSy/R3RnUSxnI6gdpN2dOKK4cfndQCMT/4JzvReOAS7EI
h8a0sEkWxirhqhfDyMmWCv/YDC40cVAXgz/ACv3a1jcwqOOmXziqIci/6B6gtc2OYpWAUSe9LLs/
5osgMqWkO7aTlwrZS4o2K1eFZUHvfAU716WbrSxvki4z/Npk6tGR9+p6pgbvszJgJy9A6ZRPVDJr
n6Ry7x2MC2ZCmftiO3QowOyaffoiZ/YKfOW++K00HPraa9x8vfOnhDv5NwtDGZC/MGGxjSEF93Ts
spoCdeJfWExikQW6eFxzQtDjvLme3s7LNkswIAm8afrQkAQhTauWhBdf/TtXTb4a4ddFmUAam+AG
dTphOni9gapN0Nrf0PkWit9jcVVDQ+7+qmGmrmaSNiWslixGFnpYCTNtYT9CbFk6tzhylL5TWqAM
vtV1gCNew79Yu9CrmvcYiY1WpTf6OB7Q/ZP2qeId7vWn9z5QBm3Mr40cj5NZQyFzT9Ij6rudIxsr
UN4tvcnqFv/OWR7ql5dwpvho2PvgQJnnvHMzEe4ACKMQlVu6SzxPJ50o1wGrPvrniiit4D9gu7h9
jipk3qZHGodK5RtEQZXCgsVfm03BlX0s+MRjIEP/FdPK1PrAhgkzj3Bp4r2n2tDoXyjec2HInxF9
5eZhoK1H3AgArY11hHr7ijJirceedYYr1Gkbg28MALCRUeIye1nrA+6pIQy6aOpaqEsq2Ls9Fvg9
i0UXYz6PpVNOcaRkcdcbH6hBMFTm2r4Si9AcoZWZFL+XRD1/MOvUezhgV6aCPEghqqD/OFTVBHvd
w+G1thcQtV9xz3UxaEhFtxhQiiF+M7YN84bvilvEgBr7ZssyohMljuiGP6OFH7qIwr8wYBj2VxLl
vNzrf24XFXuTer65ZOdM5RS633sK4+QZarkDFfh3ASmVmumQqBpJJETFgS3z5rRr7228xINxXMmz
rPQw0Gf5IIFFzdPn+P8k3D6YQZuZkAGDzPZgZ07/TkL4dEORHdmThisJqhsMWhQQZEPtA6K08bEB
40PSE3fFMuxURK9esIBYGEw8DxNhnSRdSht23IoQDhkTOh8fw/+BLfy+0LsaFew2CQG3NC7lGP0f
/6pk5zuMS/49xbWdIIWiuSYapGeq3WkVBbeuVRFy7OY5IYIPgDFGCJbyAYNLJc75+YjktE3mokyS
q02wpMMjFiVmw+bJ8/8Z9AaHgSc2ywHi25GFiJydFxgj+LOATHnXiYGcpzJ9VEso5E29RNgzU8kB
5W/T0t/G8bCu6FSF3N+UzblbFUjVx7MQPqfS31mH1kj8Ov36XlHw9GsB6zNs3fO0ngECEM1ZCGRN
IF1im2bVN8+BEk8R9J3gMiSDkbUxeU18tuTdu4WD4EZ+OvpENCA6Hne8n1zzHd19W8Own5nogBRk
5/g4ENlRMzFlmvUSzctgCWnw0Le7FEpmhuQWmmpcn6zvEZ98pbjxwhbQHIIE3mfGYLJq1KVXOFxy
AojO+QtI5Bv1p7npDYZMABvR240mrsCsQPG0g+Vc7tbxVEEHQ8m33Dc2tPl92wbz3anLKI0+4AFY
CWJS6jDR3bcvpm0nNBplq1mC+haH71giA+UkNWIb9AJhTtdk++9SC8JatgGtIg48rKrGw9bDzJtD
cCJtn93cCaLRi2MhIlY3K7fOYRui23OzAMpg3Q0mIsQ7cYDrl9e2OZP3yUhqE90itVB6ALR/NQK4
Sz3RjspqPmMQdq/GaZ6K2lC1jSIDUcRr93N2vHN+oJU6bWKEstD+p6KqiiM/vdiUoYLu+qfz3yzS
U7s3SbRfKwv77TBgWLmEomxDwBcIX1v8I5CpyRmx/99/YnXvLG7Lb23UBpp55lVzlcIUHXppW7ZG
tSva1A5fHvqDb6msNGZ8iaP4FyatZn7C56BeEa16NQBKlXIgpbGK+AiJRmBiUb1bq528UqXz5LsC
HHK+xK5Mztv+i/4vLo7U10FDmIpKyrcLxrCxeV+Dosklhv84dGfXpc5t0i13BqPm5xqo6QHVpAWe
FEEaqulgYF7rRBmTnosgxf9xa42Yul3CtW2jbVWtnr58BwgBXlSqTJHYgcD1qzTvk4fcB2LV5+Zc
yGQw4v7TbBL96NKIb0qNKUOV4fj7LbWjSARFfZ3foOfUnwyh7ioLGMaod8+5YwcSHNo/4BRK2T1r
e34pFg+bXNczQxMkeqadwXnEIpXgX9AIsNylUs5OElk2VwnVWcd61Kc47V/LHtRuHL/JAQh3FXRP
o+dMn4p3txV2VeeD/VJ4N3IBGOj/d/ishQQE/kU24DjYA+h3SEHLRaz7FJe11qg0JRaYnZRV4bf3
bY/1+jLbjWrPFK6Ys+gDFPy4pWIwp6ixQuuaicYgUG15c6cmNFXw6Oc5dPb5sWaIh/j6Bm5a7rBQ
cgvXzzSqnNGPkLV/hAx0TxtYCuOv25VR/q1PWEFpsQ/Jpn3m6dol+lB75Qj98JHGILYWeCt6cG8Y
phVJHh54bnso6DiUFtuG5f3aAJlJ+I4XL/aLhJWOUammQH4cEe7CXpSq+Qoh4hvNBrMhKl6lv7/c
PQ4z7fHD259Jv7CoNJgZ8FFs6ND+8tg8MHfl4djX8iSC9a3Bx49KP/kdWOIY+z5MJjNhTvV6RAeN
lI+OgXUpDPmHEtO5iH2BUJIMvwrBaKB/7XHcxfIvDos+9Bed7cHlZ7+4H2CiCzX5jbeOsd67Y67C
LpsDG/YcV3h3oKXdv+Te3wVwVLcXP1sJ3zgjYqJeyoIiCdY38IkBIJsuaGo1q0ijy7eWLhoqvjIY
2UfRLJ/9ZJLU/myDNY0X5IB1lLzLLKtNASHF7yiTy8QNiBFXzeOp9RMfXB5oPCns2zTDpXhdNU10
WSJLgdknmsSRJjbs/67LIvDPbNY6+6a1AVdlqaeLq61utf6Y7i9IG5MaAFAdaU/hjdk6blI7Zt1L
Zm5Bn2XIvNCtpdkBa3Cr5lyirOZO5Q+2ugqjUkErUNIgJuCAYgQO01zzPJwrOeH3tU8KazIdwxZp
q+zW9IEgcA2eXyOPz/5Ztm5zwVjQwb2GTvTqrOZ4D/l1iTCiAA21B55vYdOC+X2dQpAM8vPm6517
HNT6/unlMx7dPGRVM3OywOslfEIpAFjmeW6oV/JLlza1l1g+o9LqAkX7odEZ/6xC1EMspDuq/iEb
6owuI4A3XMgjjdWyiI+ip2f664hveBEf8c4gb92sNJvU2kfe3jSCtJVJkcnendGGaJIODWqSa+d9
LGf+udCMtP719JVbJPguK0DycpUdVN4d/ZYlBILE6fNHx4O4vMOmWqh1YddVmb4xaqK1AdbP968/
eBEUg5y7LjVy1g6v0KUSrMlDMSQUblEY5mGrFTHVAlK/FdSpYgUFh6Q+HVMSrJzcRd/7Is92IOe4
rbAFRobYes9iFw7ofILlBoQ2wiy6Y77t3+mmNmKLlZFYVUiWoZGfs5Y3QeMnzZPg0nM1vbxbG4uB
FvJeRwYLbozNwdNOigQMw8FUAT9R/rHS3mCfuDZ4CDPRc6k3uio8sOneaKPc6pWKLve/iPYgXaQa
ktz07iCFdtAD27YY1MIQTGjaZ/FkHgSzPKkdW7hpaxSBXM8DEbjDbGNO9ZQQyV3+TQoFsGeCTdT7
DKVbbtdr0jl6xU/0YjrVT6Y5QBY0ORn0ZxtPV8iPMravTgol0Aaq6mVbS6Bu96sh2w9iVGEJVPty
rGFNimggB4MFkKlyrmb7ofKcbv5gyuBX+RoMlq9tPbovVm5HFAJgZFQtonGLMoSan3ghbgkrVBLm
491HSAzDPFqi7PnN7STHme/7Af9xYI3/VZ77nGD4LELum9wDN+3eSXURvAzwvQtchYk3YNFpotWd
cqyN0+YQowDGzT5zKsib6tOzh4HycTPjC0BUDJSLSIom5PXTm/w7GrOt8AcdrfPjGZHURr3Ni+8K
8i1dWpl8JxNY8XHc9r8cpPTgl48QjjPs7ynQ3Duydc8yXP/4lYjrerzhgYdhtxuAGBVzj7xtMNV2
rsHcgSzYqBsc5+6APajmrdkvHTUHi5RmRD2uHkZojkHyrsOLJJkzmsYe8yv7XFYW57X6qmpv24Cv
fyHeE8KxRL+jO2JS/o5NeJy7dXoYpqLoFvJsvxJCNBLcZa11UjrnwQOlhRZxgbXdNqyoP/4DGdTG
wUACd1c4Lz5vqwPc7NT/txgIKEAyqPDK7cE0fUfqzWw4ODJKPTJdfSAS4NxNjyolf0jiC9IRZfqS
EyYMtKf4B5UC5bSB580bI4TjpprI3QYcKfexkOI195H+B4YB66TCLIhgkBpl/QOU8RjWaNyQF9pa
+3OEYzbgwZUD1Jrw4hDTBUTRg7Kal1nsZ5io/I9p96qeR86nBh/BceUdvMtez4/50Wiy6mnYh/1N
QO4i85LJtIPwc5ED5hf7DGNFm9aFijEtIR4Xk/HP5dT7E+TABtYSo6XHCZPV+zDJLtf7VPNi2/6e
xW397hyUF0dxu7v1mtpvhjmrYReipkTv+TlLWUUeeqpSOgf0sDkum1hp+7Hvu9bExL5opWgtfYaN
SK4q8fKydAjsWQN3534ZmojC7he2+zLIQjDJQymPfx8Ep5CLa0tjwj1/pYaP9Hkp64DXZKFSwz5N
+UPyq3U+RknyhOCYXENJKmRTEtNzMrNX7NpJ24Akoa3NKe2GdCTR5zX1Bqh2xLSoA9j66Mn87TPt
pG4a93F3vFMf80Nzy42ANVrj1gBhtnV6XDYASM+Aq3iWBzGC/ecOJ8DapKSeCQTxGeitdeLiItqE
S1BDbHxJLHjFfmt3r87bY/IweDCIbEIbRfd35ly3P6XwNAAqp3vfzYy73c3ctIRo3Xlmp1IN0tq4
BrK/fgm7bAdV0EuYs8qkpRCQqnk3w35vvgbJ7UrgMc/LIY0u4c/XFUGmbwPWQqP12BeFlxw5Xp8G
5F7lXLo1FVjhRnJgr+E0Su5fDjacROpVTGWRxY17qSOuWmEuz5Olrg+VJJZ22Vb6fH3kOFRXTgtR
n5tBa6JSmI9zUtGrPl3GQNfEPEcaDvoKYT065TXXtovJKX5xq+3Rbe7kXZJhgt34oXjAAmVzTZ8d
EXrr+V626+B0qBVOsFKY+ATc73Gwf6YHcbWaMvDhZGI1J54it0cIIddNm5nP3w5GvvYp+xcvs+To
lUdLp/Nwn1huVdghJuCwxf6eiWqwf/8F4J4l9WTiPfD/7yo7jdiivFhHetV9aspBk7F1qy2K3sku
y51audmNLfe6k/mXjx/Icgd+hf2ICNzZ+vNUn5aFehg7te/ima5kUR/5pyY7t4rqwfbB8fPb8MZ6
WnjE/qLOBtBsAwpZD04cCQ0zQgvazhh8poEkIpe4nMyXiKDwtSEzv+xaOj9Q5rDNOI24BaEnTUrZ
o+HGxl7lMuu/qq3SCymBg1iCYq1X+1cE6ZjLiSk+exXrqpVl688xwHreQeDPtTmuji7u5/WBc6D+
eUziU1XiNhKzzLX79+YM3kxuHyNhxfSKV+RmwrFK3kCZNldLdM6dt0GakqbYcfSYHEJRP5a61+vy
xxKciwrER34FArGS2chHiWSdcfj9pCuD1+cotyLBsBaEwLwJbbRTvOvED3wrnIitJMUoaCYIkOwB
tTEZxHCegXygFhNl8LfSkH3Ybn0AoO3zlofs0i1fUSiDLNOrNgnGuQoFwjiCf5llM+XktDGJNVtv
9yvN10MxwCcIaMaKmRh+iGEZDJvOlKej5ibesxhZpBefgnvPSNVjTcVHD5avtg0ZTVxGYMYqi+yE
tDPvK6WMkvSwhc636pITwxBBeVwUzcFB1e0fScxHSK+EXXZ6UI1hen02orasHGLCd96Cp/lTnExD
TgmBMSMJWZCyG4UWiMhDL9vqU+hVJ3dkWzP+Laia0kf+gdw1Zit9Kvum3iTUDgzRmNsP1uOVhujw
9f/E5y8cywiOXokEk5L+kPAPZWg5/ihpVJWG4im7q6RkyPSWNlhUTKQDgSDeX5VvPJfhkTe9ie8N
d4fc53y61U5QACigTgkOfM7+V6/r1bWUtTLLRY/cLFTU8NlEXLOr4SwkiwoKFrM+ReTjF4tpjSCX
F2rEjVxyTGCJIGV5vNHVteHOeDk8YDunBTtjAd5Eo240IK1+rfd47FimLeTyVzusYyHBh7qcNKCu
x2/V6aDghQWndFfecJAS9Rb1xFumpNa+wn8pcy1F/X7xmeKefNuf28fGRJzQeplehqAmjJyQ6bEe
2PRLxJ7cdnZHQ9RHGxOEf3oczJZP6orMySD3CtDM2Zm9V9tw+gLtmhWF1VuTc5fTmUzljjBgwAjK
MiAvlGPN7noHI2eqaVo0AjImeHNbUPIwm3PhX0Tb0AAchOYWkGxhoBPKWAhnhYC5O2UCSPRAJ5/a
yo0wtdu/OZCzTKb7bArWgZRCqeVRH1/57PDcBn+9ccJjCrw6CqAVxOc0IB1JSrPGDvYNuyojGwiO
0Jn1CljWaBS+F6w0bZOZ7ivpA1cEmvhWBLQLVIGs90O2UJehbLrqlS/m62dBLTbqZICWucUcEeeI
dIfxarvqv4MqSudVPGtJOQJX3QY+fwMkUqJjieeZ+hue/HsjWHHi78Bzo9sCbGXJjIbNwSTMAhvq
7alW06KCr7whFsbZtr33UM4eyyM4qon6U7spm0RyvHjTPdyDRbS88K4vtapIokSjYn5YhdQ7gibF
q2riYhQRD8rntRAfIQnPQ15eG04dbdn22qjTGLp2iCIQm8dPlSewvvOT/9AXyPTj82GtctORzs5F
mWQ2OCMdfrpkqPhGbqSDaZcekcZ3sgsT2ANIv4Rw/1qOPrBz1cbm5ZsLINLsaI0JVcQuGb5iGkXr
zWEErEZ6npVIOsj3NOaWNDN5KGVUuokAc3BvZXMogTB9HhoabKPWnCEl9pHFj+LHRFXLo33cQVRH
4aqxBl9+q8HeEYGsSzsiIegG2sUEYBwju0dWy94g1nxPMcdNd5CC3VsTbnsrEVyB1Bg62NIY2VTF
zbR0M4eCYlLOf4Ld9fCZF5EelYtsooYF8Hg6HCIBS8OqRuYgo/beo3I2HBAjUQL30iqDeRIgKNkL
8yQ0KAaPu1/prhvFiQVPC8B1Kslk2LN85jb6E8hTPWRRSSAiu/aBbmrISRiNvxDXJCaTNDUn4Q0l
dkSDwL2sqqhbY3qXbiG8uPuU6oZpxhfV0LhaEp/3f4q+VG2lh90Wlq9LCpucwHDwCuaSBnW5EeqM
uoF32rXYexG/3oqlTmh8UXSCryZnhCwRo9MtHHsY+hvoaKuDmWaVy8QQWTLsINJFEP/6wbk2VBkd
GB2700d/q40EKUDcn2xNdhxCcVo5oWNcSFhgcq7gFAn9eMeIL5d+7gAZWnpyOBnf0q/oiXQS4Sxu
U89+IQGde2ZBfSIvOBXtun8ADb2d9Rw0ZqZTmGGOU3y7c4CARhTSH0mkQ9xOFF8rV7R3NIh/e7nN
+xFcgl1IPYSv8u0023wupFooEqfNL8BxtTYsoDhzS8ciYpk9wr9TKylSWaBNY1Yigmro/Kd0VpEG
q7EO8Aj167uDBscCnvpiBfTJv2YnPohz1zYB+a1SeJ1TYUHMV59rh9i0sVp9nuUAWXhk4L+Mjspl
+VyPPzu5efPR6M++Y178OgLFzGseZA45ft/hKRKsehWeP+dwqwtugN8gLFx6E20TBOMaJV8qwenl
6bxAyKqTEzZbnnDYAYyOaCQGbLvdxmth4qzWZm4MT5CV09I0jHLz7sgBwVotECEoYX2sxSkUi09Y
u6q5/oNDL0407cvNaORjalWbWqRQSIqLm8PJ5K+Bj8yy1qEJuTYSI1Ndql2jlGpZKgfl5Kd7ph0V
YGf/mgfyopoXOdicYWJfu9y2RA7IGdRhzoCEgKpIAphv66OHDPTzJmLxlsZxQgHCsrby8oHnryD+
SV/4AegEb6jfdFljZIAI/cQvOb55mJ5MZusGdn5BNX74/Inl1tOtNjxzM+4T0u7h4jQKfAEm2zCu
4rGVbPMnU5n5kyD7eYpLKvB/5DSjaCbvYXxK/3NmrJG/GlCtuxujSvS11FK/mL0gY0Nu4vM6Emez
0dPLveYAvmV0lvJOVfANwyCH0n2BCZMR52jomlenDnwNtt9kqMWFc+5sbli+/TLnD1hlSPA6MFIa
WVk6qZJLgaqILU9iiLIsWzedc/pUXpkmZTkquiXSzuxYUqwpfd+HvQr+x45JmgFIp+qlMJkjpCmS
waJ6jv3xX+5yQvzyBpkQPJyuowJ2sAugbHZc2sxPdFVKIqE6ut7ZhEgBBHYN/m3T20sVKCT6MCJJ
ulLd66qdCMcB2NK/pjQIZG7QSKq/BehH4Ynef+K9n2WbRcHAyOO1suxQf6JMkGqU+9XSuDd5G7uz
OJLgd/6VuDhBrUie5boEb1tvF0Il1ndV5qsoLJsZqz6lKpUYiDaMONP3WhOMtEzEtYJ57gLQdt/r
toH/YOhwxydKTzdypYlPWuXelqW4sNo2hNhpbsB47558WPJYdfsZLOg6jsdwOzbxmyo3aFHi/0hR
NrT+8+Nw722D3aAC906LVUKNTRgjh+J9yCPc4SMQFzD5ro0rvVtlb1Jft4eXBA3rnz5wAYsSQHbf
p+DbhNLKKEov4lO595ntsoG3YOWKU+F/aarRgWU2TiOeZ4kx9s8pwME/dvHzELqtCprO9GWe3cy9
PSXSDe/wHfkm5AbIurCX3zB4UstCzHLX6uZqGfBF/oTdF0/iOv2IIZKCXJJUFFvgbaKPzlyaPfSy
oRSVBbGhnPL1b4PnYFKMzjGa/4Uj5QBCqXJ4Yd9pBCR9nNscTukqGIyviu0Y6V+whAvwz4mdZXkZ
bNWuxXPwFF2qpWxDMewl9CIJ44i9xHOwNSiaQSEeMmdYoU2AeoQ4qX8aB1mXRH1KNx2lkMGD8BFZ
jkdy4Klbu6YXoxVJO5YoPQqtDP7wUQgx3EHMpHsABHLDSU1tkjk63Jx8NICGukRXOTKW2Pdf0woW
20GGpZu4yYLXl3ngXor3UJQeg76WfbFebLDYSsFfskM187QzS3wbk3ruRUqYoG1BYmKXAp4YDts3
tCm94ujPDZmqVxH8axW10RJZI+ChDKZpv9ZndGIUw9yZEcJxE3cBbzvgHoUQ5A8KJHaBNPjzQPT7
evl79iTqlfQ4fWW6FL69fOmijJYBj7X3tkTt83pn53s1QiJuZ3P+HGarotXGGQuo3+2/T2zcmptM
z2QmgmjVbsb6wm4pnpkUWldXuWlxuKeBOjKeJwehQdkMCT35DLTgFcptrkhQ7akhnScsnhbdGGMA
qyBkNYGjNmfpylrgZ56WCOLDsvyjnFhImGhgLCOLBsOpwaQMGlWjQp2XukWEkV8y7U7RnACIA7au
xxYTj8S/IertDnRlpNKuFecR+XSv7dRg11EzpIh8sdn4JnNkgoyz39uExznWF74dUZHRD9pINh2W
rzAP2xSfWZvKwZ6xfLOqEau7xWIwCAXh+Sdi1ay3lN3PF134q4ELpMA2D7hUniikTEhGyyjNLWb5
0S7sm/1XJNFpjR14tzuQlp724qDG/IbjoYayNRtJu+/wctSNChuUL2LARTzhT79jwRApCAC5hvIK
ye/t7lU8GfhSm9cY0EKiHe9He5geCj/MJTiAnCcr5K//D8E/P+Po8f2o51TATSILpk+Go8aTBRB4
FR1QzaoPZZQmh29DUCuIVWb3ZUjTtGH0jTh7rVpCGn0l1ohBArX37+SOm4oe0E1Fs/MuocN34lNe
A2i1/UBRwXOVg+EWcF2i790EMLjojn+9Zymx72jAHdtXNM6DQSqN9Th74fBT5oFlMtSz9wLPfYd0
O3e58jTf1JtVgTg9UMTpF1OQ3w6DRKjenY8T1fv8Q7h+XJeARv5eW0ApwktFx7NO8UZgu+Lcw3lR
X5PJFrESLONW+GatOqHao54r43YA5FISPzBnL9Xhw1oF2QxmgNLRDHEaDon2XZi8CM96cVbLVdma
ATOz4Nq9lFom/8BrP8h1vsJa97l03TpCbeOxu16Tbffr4eZpd8S0PgWExtm/nlQB2wfyMb5aECFA
kjlNMXSZiir0xu6esUJiRYlGn0OI40an3WNoUx3w5Gtfm1WrnDXaKcxnJtsCuXjqx4wvXRLlleM8
syT27zgzVapFU7+7H5Br8QLKimAY24G28rCSk3/aekhKZSEHDobDKn/B6oQYiAAHS3URH0hISyVn
tqBlpvqcij7dlq0JhHhnRm6/6z+9tnZOOEfAldAqF2tO5VfCKloCiWIdxc3tnaJro3SUlY+StmmT
BDmWk0Yq8Phgf+3eaY24ESDJvhbjSsOpEeG4qZ4Wz0sceElenVquH+tKyxnehffujI9ixvnn1EO4
pdAKStH0OHV1GRyD4KY6M2i9CZby1Yvcwo2BQxYbxeQN0Aw+Kv9pnfIdfAQZAubS+MlJEYXArP/Z
Ka7meod1EYVgz+T294j9qNbgTg59+Qpryyvj7cG1t+sWEg0CgPM6j1FrhDXHqg9j9fercWbsYe/O
z31TcJ+FNU54KiMHMLm5YZ3vh0Et38lFprJFvllUK5bCJHh5XkuA3vFp2Z5/6NU18EL+B0ir3FIB
LLAV1MxaYEjACjU5emLI2M/9AOhJGhe/+iKU7as7HCkaAOokiBb2Y7ExLXv+rw2Sfdk4mbdM226T
ZjtBU2bh2RjVU4d2t4KtEHwY1AQDYBznMlsknciaqDBjf4OIJLLWKcvnHo2eNfa44NjDBICifvSs
2wlPrp2bsoO7ghpa+jTeLGDkbDFo6anqNmz91gKxYv0a7KjlCtv/o0q/LX4Np8qcirPe8b/EOCI/
k5+m+uOYCjVzps1Yi55X74lPnPrmh2mMNI6phi3OVo4fHvdPrc1L1R93X+H78EWYIGtPvAdN0e+y
rteD6pwoNLFBXLklJ64W3JDtkXBqZbrO3xheyBS8F6C7MsA6wbJrSwDEIC2mFbVnXvF+2hPDuUOE
Wb7VyRjL8SJ9D978cZRQ7MY015hUmzliYV1bvj3Kj6idgwNcCm62x8DzbhCYMeng47syk63lZWdI
a6l56fLKZ5FlVkMZOCXh7OLhz0BrcdvIEGmiHVXkppRPBed0cYz8buNKUfMPC1hTJjwNRMxAWCtU
E4C/L9bmJ3XhjhZiiWYI91XhPpCq+o3nrCCHPvjDbfgkrUP3PxPiflfYwEtTI4HCXTpc4ubWIKEo
Pb4FWP61gXmeNPaoFpmCqK45rg8LDP7w3AVoHX3JH0QlRKuQQJ8a301/CQTzIhMJ16CXx+FNwaRP
9e7m4OSWjWX+HaxQ9+MlYZ+3YRFHhpNHK65dBex4nbuR/09vahc1Ctp0tYDD9C+QPZknxQW1ouBB
AgHfipp1qwBfT/59LRUt9XarBV3Ra/hqU2+uazrYquEuh4Bv1P6F8/mopNhFacpU2acsk0ooy8yg
KXgIy3C2FJOFalv5QiLoPNNVWhoZeSmpooAt+tGUxz4YOnXudZGVe4RDaKBzKIiOgJbYyAXqDr9H
Lv+wPuIKWfqQVN8OMY49QssddqCJppGqKgl+wvQOAJU9arpeAqDqEwZr5vQGn/EOzNT8IvEsRRty
q+uCOn8l1N7HmmwZaypYXAWXzcf4YJTb+/vd9qkhUOIW1KzGHvPwa8hpWM3ZjJtvbCkCeRpLBXt4
0p48kKol9DQREyjGNx0KW4xRxLJESjFsoYUnNi7G/CVUWasbQs4Y9nyEw+vwrpDiRvgs+n1/IN2/
4Y3VdByQi4/Q37X+f+t8/8GimOGflhcq7H3pASa6Ta3HdG3zJgdu/UShkj2coKu9NQ1+BW0ZqZEV
MJdljuw1jWieAjMq3eCOHcJqO4d7vxE9LUiQm6d26DccKNRGmEU+zS6/GnsPnbwckZdGw6+sgC1r
E9h0HNbdjV1jRL2ETdTGSPpBC1gk1OXzXEn25EQGwBp8Dkt9V06jQTJoyllSeQFjveMQSJMYk2Db
88bwpnpnpDhTnJ+XKxJ7vE3tThKCYbbfGGj/RyrmrWmFQX/wgDNJgTnajCTkUTcxJ4cGUfZwbRbq
7tFYq+FC43PEaHjojd8DBaMu3sFsNm8jBHdXlDEqK2XCzFCZPH0YNcZQElvdl1WQ3mhuWAm8qIpw
MuJMYcMmAeSHDwGS14BkeYcDhCdkKk3dRQET/flmsR5MNk/FUq/j0yE0HFO0qcaaXdY2W0tVOyWl
L+ReYs5wLHAUdi40KH+w3LSGA+ajgIbU6hQm2YSSgZeqslemhlX9d6Q8uFcBNA1iwPjU4l/0/E3c
phwulwhDL06vX5dJ7QwPyYx3CjNMUKli2dYpmmOAWglo8+L/nhlQ+BuOeyIQ1Up2dBKk/D2ciH3D
l3bnpz6BT70yJt4VMQEVcK1eYsYB+8U6Rs8i4tuheoIeKBgDZuPiEkLpMvREjgLIVEFqOBZTJ1Au
tkc9Se2Dbg1iBPdXVyI5QyKxw49BvCac432sgjs4Gj3WY1k/1jGPehA/dqw1p9HjaA/oqxyRNOuk
KYrhVQ0SoZPice8MNVulRquk+vgYzsojlCsuMrOkcHaHBQ0Nm0hF8qUrrSt7ytwKAa9pAfJxRd73
QEaGjYYYgZ91DIOHzb32ztigAnpVxQVrOyKYuFEhk/EQLQIoY3zMIGgG2qCasm2+8uBa352smLQn
91jidoiI9XUuo05F324zoJ59kBbFV8ZoE2HY0BRSrdKx9XF+3+TAmZMGB2T9ovfDTdkcLhPzzx05
wTqxuP3U9JArC92rbfLAoc76VnxV6jqjrdtkkwl7F5nHUV/j/j2zA0LBS6nGp6AL/IKML7MJ/0WN
maBYMIMeantDo2nhJJTxWi1S3IWp2PaqdwpCOOYy1M5u8oABuXf3r1w9oOzLej4kgeWoAz+zgfIW
rjJnuSxPEfCG8WRwHFdaDmAE/vgLoYoGlmVB5mQDGsX3BlVp178R4J/XStVKUTH8IEbINhvvAiWP
DuUUyeT1q8JAKsNNi4WBeIsFlWDZcAg1PyfqrXAGOnxdfVGTsdrBwT9hWzVgYEGh9npTGyxn5Bv5
yvncC09ai8BP8rAym2q0BgZD7Sm9U4TeK4BNot/NaTQJ3SIlrNziGrXyx1aaS8LK/gWtEXoVrwSz
XZx/5KXg0erI1P3ZvdDSZQHO6uQe724zhiU1q9YoNfhABhIxcwIS/ftYk56ymy2Q4KFdu4hWwC7A
pTjZEbIFu+P1VEJOCaX9ZVc+JYyQiePkFz2bNRlV8Ub1VYVF+69FHMjQXJ18gyWTCDf6V5r8wZjN
y3aNWDlND6JSjQ62cJxTHnxpTOO6gKO773we3HUIreoWI5CZxHaBnS2cZat77DYHC1zB4KW7WxUm
ivdSQYRNyLavqfpzLvRnxpC84zxlFLFbTkzmGJ7vGb1l4DdHdgstX6b5rEdfSR3Ij5m3ZD8kUuzz
522CiZkoEO8iEOziKLpLc+U9lr7/JZ8JtYio3cAe2+5ib+GFBtPLBykjDq4q2Y633lG1ajoVRWj+
B5btHRkLIliweS3RWGUIDTJdP/huHwcNeUHWfKSZDYqiv6Sa6vf0jca0aQAZTUtBxxHyG2ex415h
Vhvlk1I4UtsnxQnxG0cvSzSWrUiPnkAfyHmwQAJOwvpflOyGzKrq6NpPVP//ILY7vwpTAbSbGqPP
0UAlCJvVvD1hEP6Pq18DZwUX4rs2ttc3xE+rafWRtN9PyErqNlZcdwKfuP9poj9uQeGJzbLnUSmF
vXRHv1Zpk+YUs2b32k4zioqMI+g0ukRvIe1OA678MPNfREggxvNtx+nwn7Aj5UWvJ8qhz8DV0BsF
NtGWIGWgdBC+zIJav+bNniXTR+qFhobazLls+EGeczrUZJNEwBmijTQ+rMDERYpHkwXkA4kKYT7X
HHNmAMFZRQmvWEpsU9tiUTCIFz6HClB01Z7ksPXDvg8pzqYRH+uxNaMBAaxGeHNvGYULnzLHZh1V
9h72stAqoiKAxFZqAdIy9HmcMgVzaQBY+wXPR59rD/NU98E7/FiZwHoCBK6Fw2HlNnkme864IoGc
nSh+sY6UaPo1lMsj78Z6yAWBM/v29TeL8rD6FMUU5sogzFSfnr6drMbBZ+eY+iCbb7hmwNS8XU3V
CGTK2YMvf/qX+oLl67PKAN0TgbuupKoMes23s+xiRDwkkpmL0jKlTFxLvexRZpTNqIzSuWOawAvX
fP8o9AZs53SGSRGeXgFid6B5t7srtRs0UQksFqouuT5Om+uW2tqc+SfGaN2sa8RnPhj7zh/Lpp7l
S1yvOGeQ5BzrWrJKU6cYjkUR389yTUsmqwGimYicaNl85j9GBLJbHIgTxXUqZfdaP/QiOZ+RdhG4
QjY3TM/5Q8UwnT2QJ/M+H+6nCT5vt8pmUlK/7iSs7FoTsACjbdpJ/dSZZ3NjAMi5WFBv1h/G/Pek
6lMlATkTMsT9wpeWRkvw1470JDqw+p9ESsznXnxA8RYHqWopM6d/RwOXGdd91Hy4r49uN1HHdw7c
FwCiSZpduJWgmqYtdbl3kg72C7nIVyqPpdz0m+/MSGSj4VqfuKRwhp38WqYeUHQmncTtkpizTJrm
+qZS3NX6klIuOQtF6aPBm6IIMgYBt0S9ZtUxV4iLzHxsg023NV6Uo1BaTikXue+rVK4CMBxx1Zv5
s/+QAyWEJI49iFyy817jIVdbtGs1jAnrq8fDSJUUd1znxkoxYJY/+7BdgbpzzwLcANwhyKwjpz8R
I9LHP7eIgi43qviBhKRJ2FFzXyhzEoDSUdfdNJnP6ZNFby4Q0orod1v0bEPnmWPm1W1sNuZQp7bP
karj/nFkjvP859y069rOyWhVgLdhSuvyAwt04VmwBVpTY7tmXoTJ0DiZ/lgK0oksfbzhKhYLBNCW
X0W1mFWoQDi4zqqrQnCt8a7dywdPGiQlpiq/GLovSIkEzFRQCUN2LMEQpLDrUPDWgAZrQGqiEDsz
djCrwjG4LSGjMhtJJTlHK4KErRiKT6gKzf029qgXcvkmZm2OFCJkDJWGp54De2NsTVy3zMaWwe1L
oBoFXc90S40LW353Pzo7N74uWHyyK3IQRWGDfW2Op69ShyMzkkrQUQaCdwcyAURvGLUv2rEt7/7E
9u/x1jqLfALfLyZmRCBVLmtKpN5Huu6Ony+dlo5OYdo79hPosKN2Cbkb3cxAieJp/QN1QTPMG7yk
EsFbSHtOTwj+dbQyU2CjAQFU9KCfIDmk0HuMAlE43rImxEDOOAoFK6xfjibl4gip3hyM62Qk3yyK
OuPSf0gq1ahkDxtRPThNKXzx4lBh6dkvmxM0Z/1S7nsz+s6mlB8V9rNYXbGje+epTlQCnW+5m8lr
6WXouPi867IS/kLDPtzT5zSuvNP2ybCgoJx7K/odt8pKTUe5PTg0127S9tOHQvbDB7rBpVco0g/j
lmlKsoTVerq/SlO8KkcT/K+dEE6bOUtR0MYzA/HvqOR1lh79VS4XMqd+cXfZ4mxSlz23yluFY6Hm
HP1H7d0U4heetRTCCU8lGxmRWchVXH9iSesUSpGfBvb3o6Obvj4Ejm5nep1J9aRwKFtfGpKR2rTa
/kPKycezumtvORT9OUtjpLjdrt3vpitV3sAE6VliQsqHDvEjG5MCpEvRYL9UxjNyz+mxgYLhj+YS
Yut+jHREa+syZ/wTz6IMPQ1zZJfEE/xRVYo5eSzn8sfQw8PNnXR74+DUMPfrC95XIKdKqfkR+Xtm
d009HjoH0wrk9oVRLIHHEVlJDMhHSLbMboebVBYgB8frdII67cym8IVW1v7umJtDsQqWDIAqorH9
GShxN/yt+yBPbZczqpvwHzt5Pbvi05HS3SPMNy8FXaphgJVH6EgghdAhBEHpCQwsdQPvwdSyz/RN
IMzqvV9n6mndZUP7gSaP5OLIPd3/xawNdV1yQtZ+QjZbWt3nPZzK/duwuhvMU2Gfx7H/y8lmzRwW
I3nDwwrznUtqo+G1AfP1bnZkOzEI1KSd+/GVJ6BDBZphaJaw6SwXdizcckCFABJhF37FreXVvF/J
V1NUXjRjVRmRnOu0tJ5hNnp4y8ncdveAmtufsE9nHLL4DBFdKv2Cp4jwMD4NN4tzzIrQYI7GFNvh
CuxFxu3FDyJrrB2Cs5rvdK1jQ/JmTcHVb5AWohdtSeGxwVhp58wB+C3gPUt44mA3WvKAOGA5lp8q
AiGviSduDJQlO1Ymo/KIOwWghfeURdwx+cOTtib+/19t0RBWKWqhz1/cWUXXfmBYEET+W+O3sPkk
gvTBpsW5bzxr6aZXxh7riLaq2D/nXtlOx51rc9e41R5hfsrK3w5hO3C1oWlGc2iph6H43jwdH4WF
8kvFn1HRXB1z8WeGWfmfLkp/z2Tlb5sfFEFoEn0/HIFwgIwHEeHRsvvl77sNLFFuvlT2wsQOTWNj
9pXTjPEz26P5+0dQcbw8lV+wgT0C57QVjZ2QiczTmL6JoIFPFHrd5ch/6JAfTcdY0FBj46RpZ56g
pCQ3FQLNvAgQELoAl5kN05zoFuwPKzfrczwUS+jvV6tYURNArHGKlfZO0EGD56665e2hz3LMRlKm
zCwC1fzvqfURf9GMxB2gzcialZf6fYI4j0QtSXyt2shDUvMzxFVoy+YDaK1OfcRMzjc/n+VH9mQ3
9FAbaNmWGROWymW/q/PallJIMphcMPjuBz+617TEjy00brpslaQ6/4iiFbMKVfsmPPv8B7rrEYsD
IpGHndsbZXDCaOIYtOqHHi1fkyJMfq/aWK0nXQd5Pq9Ay+TF1gDP9glwdsDFrNHDGrSoKttw7zr5
ZOKBEc1qOYZiFEQtRPmQDr/DmBZjz4Bk8SCVAswgQb6hESUtskRbPMWG8s4YyS16hEQpiMm9chjr
Z1nRqegIHz3swHh+2e8VGRIskeT2e0oLAARdUtAWQbjJGJwGfdJOZvRiYzyA0Fr2Zg5E5vcbb6zc
i6b31Z2d9eE2NGoYlyZDEi7eKWZH57R1LGx4qvktwQH34/6vCB6IInLMBtxwxphH0L7E/WlDXAeA
GcbD/3Hf+JBoNt0nesLtQ1jvUEXPphDEIjFU6qOcYD5t4x9OaUxQk8wGO87CKnIhaWwWSCjRzhrJ
HsyEFZUY3O8b5f3p9T9gLXseA6RopXG6wfnvC+1/0m4PlVRAgYH0WlbgvkG6BP5c2mv5xuHmYGck
BwfAC2ro40MH7BNey9nlSWNTLc1rZTkCeHM86vzZ/v5yAPr9pqxBo2d6/NqKFnIgvP1Ckqw0/KKg
cW3QwNObCahey/F6VBChoE9G86zz6RWGGBMMG1N5wk87iVdJYnAQhwgUujgbW5q+M8hhRO1P3TR9
w79wBres1TRgY6FtUT1C28dRuQHZQRjlRjxY4CTnqJqWkJxhCGH4mMuFTebYSAhFsErSYXtBENGO
x7ieNEQiNEJI6yNDbtJcpbHyoSjI93GzJjSoQISXiWhU3GzMrgFePLLOQUuDRMxkWcXoPCvfi/qf
DabY2fMwPpG4jdlIdcywaymAx1seoL7jmiWicjHBCx06JrvpWQAsui54egysIt3KFGTeaW8jo8jU
lNnxoizeV4Vn3uehDNcqE9Ga561T8+v669kA7urjNGIHq5riRzL7fIuhtIJ9H43YvRjQ5S3tHqjg
rigw5EgKZ0QlO+mvBRTmLGUFhaH9bwdqSMzjRy+uHsoChvPvthib+eorF3TilqAHuVBMJ0pe6ie9
Qi+/EqNr4Mn8dPwO6ctCkkyIOfK0frRhUo9fd6btFChmAqSLP6PDUPCTwSo5Bb1voNEV/qGEsvZB
te9jZ9HXBphA+uVn8QPYX2c6PsOLZsH0cr03flhkM/mmm5npwcKZCmugkeTvEeDcP/gWFFO0wqyn
20tzzezMvEqa+bG+puVaQl6qeIhbCKmLi9BLGuFRaYN+ajsjKqgmTQunUigONj7J74ob7F0HMeor
NNjjGSxPyS8/n3xl+IK2Up/WBtaEXf+VeSRBcehK5ysg2/RwLgAW1h04wLtpoQUMhYBRkg2FEFAM
+mC71ME5IavI4jUSgOSaCGLAPR0Aa8vn2PrTQCHuILo7wT5fa/k6ecnoktwbi/KgpxI0ZILG6ZFa
f8TlytL867vG2oJiA5UGqpctpVXnEOB3RMWVEbEwzXlziAHCJfyejPT4MG/t3gqJo1GtyNu+23r1
ePmTbI19SDPzyBbKcbVkuS/bsvGvZ15vJfV5yXymqUVwhRkNxUWkNEfMb+HoCEyn09WD7mD1Am0k
uTlta/eEDSw9N4/g2ZubVmovQhaqBxoH0YgtqypZqyvkJ6NuwuXUoNOxcUrFP0pjmTW3dKZd/F8C
em279weShTWU+PComlGtcCYPQoXX4jQuz+eBSNjmNSOj/9jaPJj8JNApl/Jqio7W99Kn6TcdX77F
EXvfO4Rh908+kFnIZXX3O8EXRl4daOtG2bWCD2hPAwS7ipLQlhHey+JWKgS2bzrJQ0aO0pE/X8Ao
GqyptJCtfpbbzxBR3MgrOGBSbZyjxAf0qJ+1Rs8+UkiOkpz9WpSbjuzObTvLgcPZYkYNTwJhXhfb
tCbMaKqrPQfHVsuSTsnfpyuZDDbGSmepkxN83nUE5j+0wh5X4o2+cnfccgyNXzFtehwlYXdndXHi
dp647Yo4CLvkd9SHMezNYZa8NSMEQUWyTq4tTlZzJ9mpXt8rLNelxOsR1JtXeWPi9QEn04TJZH2B
1hmK8JqOaxZXWbgaI/vm/axjm2YR4PRo3Mg8w9Z+ee95Erv36TOJZAAkaOMEAF5jZm7sqWzOl1F/
4ve4p/EofR0VTlQ8KMwv7Dw5g8APp5+dRXjTOJ8kSAlnDlG9tdlX4DXNsAQUdREszQdzuXrWHJ0h
6ej0sSZe6JI+hOnpdz1a18c+rYn2POpIiT/2Q/Ln24T5M6FBT+ug09VvG18GGRFYTpHPxZGTTKwz
ab5hnSdgij13OpIsQSEc5clkz1CkuM56ARjGyboUNmXaOd8lrdVwL+MJqCESrgDtkAxazsO3fWPJ
DvnDVWqEtpj2qICjc2SXbZfDJNVRz7pVZe4T3RKNI1GQvPUSa3Szt71NUFKX2qbXWv5EguW2tNbQ
slJsvRyhs5KQdNv3oqGJkOse+DUEWJla+IcIrLrzbzexrWvCBVyFZuw+xnY4h6MjRvZKy3v46WA5
kr+sZjt/2S7kbjupkXjsgVvWzobCzzIPLQdn6cZHgg53swC3uh9Eiz/ki4JEHRm2e7QZytCfjZou
jSiM1d3vRAUYmUpxnbIfdjPUy3fuGUIqJ1IEow/q4uw5vCYqPf7oZfm2IRL41WAR07lUDJ9b3f6I
TKlZLdb2m2oSQ5uyef3QnCD6UT/0muIIid8HS8CBlWC6s/otZh+1S5YtJUNHp4JDqN5MkeMKxsPm
7cvcw7suw0n4XdU4Q5WMlDQ/BEaim/hTyoxvYCjl6mAr1zklYfJTJXndwPJ9EuKYPIFn0vRZHJHu
dZ8WqnTbKZQ9rPhtyI0B/npOO+jmkag4x43ZmFhooxsrN645EVOeYbQ1sy+HjsiozaOURnYwiUp0
eOv0xraZ/74ew4OKl8nAwaEeI/YnLQfm6nPpHnGfAVfUHdlXZugTvpJBHyFPkD5Ip4fC6JzfHTIR
SMzcD00VDT6CTgfpGdHpqW17sgDgTj5fWNlIZLNmDT/EtRgFbLgzQVpJ0G/01f1xH1XOMjbS8J0c
I2dc/zjo2hgv2k7f2ONkuoNroSj5l0R+lp8JB7F1aLPhvFTNMv8qIkYGwBLjQDpQNkpb9qWr1sFt
4Gv/5u4ffe+KKxvwT0DcD5KeOC55U6f2GdOph7bf5xAzAEN8Z1GpArnE7swoXepOMtqgRbZ5PlbZ
jSVUlT+E3gjZVGBz/Ga49SHIobw1292POeT+XvlW/8+hE9RazUt1Ntnh48LaMtH5V96OpYeKy1GY
BB9nSth7oy6FsxLPjaz/8mIj9gnl7QP2t7KtQpYSTYSOI11FvJJDwBmpKGHGuIpg45lvLqlPotVq
dBApTSAcToOd1vfF7+5N27l/NiAflaAer0jy8k0Ubux2Tk7H4PyKNondZKupnvfgigcawV8MZT3T
O8H9y6W7XrjSaqqeQDYiZ3gpaqqohA7tmF7DtsYVMwWosmiakDq9lO5BsFLQz8veYBp0R4CUtI4L
LEUn09qb+9cLNnlUtRgLEajRcbZ16rhEdoPLB92N4Al4s39mBGucRE+RuxWbzKVLU1T50OLxd6vR
LIMWzgd4EsJK0z/0WeLmpyeSw4Jh2XewEaBzpOh48grZZREIgcbWCyVBhDL1GHYtBzW0Bjw2WxTK
Z6XMeRm3xmrgWweOVpYls+mXJ4RbU7NIm9MQ5Y+t2CY9dPSFg9AWnDfua/aVvzccYuL8tlRD+aOw
weWVzTPeZSs9NT3giQVpzLPsxWofvVLergp9mggAscWzruXY/2lpxIhDk5aaK4KVXnZAP9ilcqp2
zLRtrq5f4+ztgH36eRFjtDG/W7ItwtyRxQ9BokDwHjMqGdEOmK/OVyhXGSWXmspjAGqsBaOqkYyE
0y5iLtcanFN2K+VCfws0iGnguHuRwt9PCqGc0fT9Tz0aABF9AXPmaKl+9rn0i33Gag3sVVVxvxa/
m6SbYiLtEuvjgvqf/OUeU3ZuIjNzVjxhXQYdzKVRdIcbr3xu5no2cBhszsF9s6IEdGW/vwLg75cV
stdjEQIFRy6bbkjsqHZLjhNyKOT3K1gM+LWPVwdOIXlnGZQTW/9cCnd4QPHfPV8H2HD7A7+Njh5l
OKdM2xXeCShqfYUNlaZor583OReX1C7AW79Ggnn9+CQOjr2pdB2gRbsE6E9jnBAPw2GllUnOMFsB
yY1nHiXbvmmE9HdEUkvd93KtdQ/en0wbsMN9UsjixTSt8fbwHuMD/dE/Mkr9j0mjS9VSLJVFFvvq
jpPRJ7busxZob4e5eIsGh1EQMalgtrgeVv3EMiKSW2qcruD90CU0s/4x9XZn+wB+rbZMmVK/OTNP
DkiwFTovCMzOziZ4uhJRSZk4So7QFR4TJ8035E9xdxJQDxgF+KkY6TLaQ8po8crrux5Dwnq2VfJ0
72WIy1N/vzPScLJkgPfNQsuDo//ICj2C6WAbbvA65dqNU5gLNSTKeXCfYpbAgE+qb3bBvJq1gq5H
Jw5b0tyaV7sOzG1v5x3nIyteqq1SwVPydHKubc1PjjL0pzlqnh6zOjDpqlVtwgvCDPZHQhqCjgzB
GUAXBkWXFRbJmakQqwfcjmuefSpxQEfpsgRntXj76zCxUvJCTSlhPfRvdNHPEAddSoKLFWKh/wFS
1tHJHu8t+XwyuChNslevU5ewhC7R5J+pp8xjtBMqo8ogAuo2VnosFFWIVYw7wKXWoep5Jn83VomP
7tDMX7R8DfeaNVA3tJX7CxLqC9cVN4xlAoToKjwk0MPUX4NvsoV4+K+hnxZg296c8lhul6R/zUS7
QGqHI2n+qycxI4RfWQUdlcOemvuz0JssCJq47IiS4d7RqQfXoVIF50IlqN8sXDPddmmaEDx3SUYv
WL8FM/yDIwfPOpKXPXNkb9PWwF5Z/HHRbjbUIJuOLMO7pTKQMCDuS9m4Vq0u1Dw/gVQYSB0HfoZj
HUBSu4psjVlExZlSIPWCHBdc4oX2LJ45CmRxtWNyw5qKO2S8vKeKF8eT3l2O0Xu/AV/Yc7VYaKxU
QMzkLzjYGmqFYlpzkD/PaXBVL7HgDbJ54IU3B4JPyvnPH/xaqCbGVnWKr47hKgpKjnRISXx7YjTC
Mx6VgooIZlvfNrNedHLDijdLevcoesLxvUtVdiaJYo687VqxJx9Quc/jvnAg7ZTrfpCkTni4mV9z
igukm2xnaVXWZVInBuGuEj6UtdmqUUkvSpl3+y1UtGwBOmAP4YUwjT9bxZ9mg+BDX58Vx8WfW+im
RhOlzaF/oUK5J+1TEglD4o58yM3thMBPlwZB/GOnA4mH9q5MhWhpYdpTAOsX2yhDrinj49FotJsA
a+0xcZxJUAHmcPrF4eUReNb6gtdS9f8eABX04+68cuw9t+/9I+YMMALy9RjNqOebIDyTb6b19gkS
KKVD7+XUbZZJ1etq+A3ZCDDjn7BsUYPa9yUH6aIfmWO1X+m2BpbBk5WT7DQv+YrGznHZH4OcIGha
qjmDTvhJ6RkDqPloLCgaeoIDOaDB4tLcSEYE+ffdPaea9Q2GlypyjjeCFpAU6mAwQqgmoTQeOF2K
sPNrIMFL8jlVselpcCaQIq4vtrRv+6OpuNX7gjfoylMOGyhMMRwXJvYKysBBWPwaiNLQSyb4IsLX
cB67/jHmUnezuuJuRXzvgsZ2aaDvfjo6yGiinmOwj0O5l4/36mt++Dw4Oy0o5C45q8RiyZlLWV26
raKk0an15tfejLMB5pz++RpEGSPK8XmV6jwPJXENlQiZg8nlJaIs8c/eGjLUkNAnuSDb+8ZcUQ6y
Q0Sk8oqbB4ovCcPPTGluaXv8hBe/Z1J/59T9QOWapsRMbjJyiQdknf1uXyVE9INkEOCDzEtvncZK
2B3C+j352anFwhD8sepAE1o89y2iUyZzf8+GHmk4u/ONUacPrSvB2AwM4oanphy0lHH2wAFZMKws
+nPipWWXCCFY/MhK+ey2zkolBdDGJL/H0qAOJCJ42gzptS2WsEnU27DNUruskVx77XMTzDOtA/wd
swxjPLmRf0+nOQRQAZpzrqM0XnFoqKx/CyFlH40mJwtzFpfbgAoPbm75bkMQbT+y0M6nrE+mC6wl
5EJlhezIvJOIOGBvcdtsyR0nVRVSGJ15XDjIWXp2vCu614Pa9ceLA2/V490h3iOFyPN+ev08DAGu
i7USNFXMa9i+dyfBFbmzrkmxGLgokUm9vI2Y2Pdd1Na4CZwBRD0s0062KcF1rw/pl1GtDySvCGFb
TqsvdKjvSQOgj9KdEzLxHNW9MJMLOnjZbVgyLR2yAANTB6LAhEv1zlq3q5d2g1giFlp6b2m4yACU
PHVOWgUAJLu4WckFPOIQQJAlLosxadPQOjre9SRURWEu5Y0AenKLhaVNzUywN3PTJnVUd3Ch6JWT
u4AE/JzIHCjpGvwI2Gmpg+Iq6AyXbqqCHqPzhjgJqaKCKMKDxmfbsq9i+HMxTWsfijCGomYNX6ar
x+uuH1ugAARswzvboPV1/xOx0xTwBhEbPkn2JtzeSqTNEYOA91G6ayp/hOGmKg8nGn8n2wzBerhN
qlcVD9EGnEFdMARdofFvgl+MX4xtGVM3wbeoqUvUAhwJIiOBJQeFFfCMbdYX7fv/CHrM6dH+rTkr
CgDy+S8cSwC8zLiQGDXsQRZ0ScOb567vNOjfY55JfKaUax7/s5M3cLEclSM7hYhTMCjPLK1xsKCX
+zDYPVUQbnTgtOyT68djZq2iM2lUIEO8tDEYJdQHY4zku4AbUCP8o4dGqM8vDV1xC2kpu9xLhq0I
fxDUsD1EGl7q99PEz+xVOprUDW74KRYj8925Ys7s06DTIMJrKgYOqc+bsBqCiBx64WHcsSXbQcNy
RfR1lnnG6ucSO0BwjEj2mNwKb1Z8ugQKZ+nZ3W1RriOzXD3IChjO19RSmRm3n95Bm581K5NXg/0I
lSS/euSD83YG/zf2pd8Mos3S6FeCabiFOMfnHd18BQLxLLyb2mVpYvNiHXTtuw8P48w7DJQ4vRfh
iW+7AlwP9J7mjzGCU2h9Mr5echspOE9N7HF+oeE3V5UkdIAaWyGyoggtYjlBtRcxLwoXkrMmFxxg
14qGDq+6KiNWPkqHGWkuTQKDRr+W/JukVrjrSPIlm7CHRWH9gIItCOHwwY6qYSfPN5TSLraJ/YZ4
Z7+d9V7cd0EFBNPJVKihlLaeK0vuRjPPqZ7BckFY4Nf1+Hans2DVN6vQ0AMNwBaGx3CBiNkyo9CD
FeUU5MnzZV953nxb7zmOOgwrLkfImEZfTETI5F+8eSCNOoFmU7NYqaz/7sYExYwK7Ry9ZjVUF5CR
zxr7NEr/28g6ffAkeK7fD+iYh081nbfEcaOVhgfztrz2ivm5NysLxvJevunMGRD3fAgj8mFAUzJN
JRPso2H54IRNtOzhnkqr129Wya0r885iz3hkgI7PDJrkPTdlzlepR8yg8qCXeglnGGGTGWP+oRKX
F+wovSzmkf/d5VbYZHnMxXDM2E1LaaxH8CmY+A90+ENj9MR8bjWiAwFkUjFTyL2jIoQUseLjyLei
mT6AzAoDyGyXzvOoCBxe/l0WgIKkNy3y4zXR9FwQB1b0IZf/Ka3sWtVXrKcHq6gKGy9EGN6YAM35
l/2f47pmkThRX14TZMW2oK5sPJz+CTerkjn+qutAu82FYwo/VvvVmU++3bp9nNkB6AgzLq38hQt5
Ji531XtyiYr0CIlslHhnTkFuclVDGLdLNuJFEevne4FfHRamnupLnHH43ksOYfmwnL0wI+ibB8BG
Abp2ND+yZMnba80VBXy2Os9RomAoyoSu5iRIoekPe4HjUx9FiNcxWIEirlFqzVnomLUBWMn61GBZ
HZq9kGG6b7vkiajX5jO1KVHDGlPsHhhlVZS9AKpGRbcMzaMgOiHxc1ZE+kCsnjoI+R9kHI6RtdBz
8HzNkx/1wjdZjsD0leOwYbbvHgxipzQTPCkuu4/qhudglyTwEWb64pd52t+YpZbllTRDq66tKFE+
Ciw/m4XH/Rd24oz9Ts+2azt1n7fK7zfeiJcLFFVxu1U2dI0wT2VKtw0Yy7srX71CSTeZZqBeRjZE
vshPEfj/tw7kM1cvKdM/sGMTBrV2P6p16CJwiejY/3Qgk3Pzy8zDCKYlmRKfDGlCOww4/GN6hwm4
dDNh0z+EhD8vyQIOEXjvEc8mAiEDKJHJyxK+qj+YTkGErw8Fu6GuvFLP4PdxIb30fLoEMiVZqDrB
sX3EcNAH5KPrtRR3EjS+YlxWwQhvabK9507YHw5EhNIUgjYQ8QXyD2FG5uXTeWkV0wJSuJdlQqIG
kE9Nu9PchNeuxKLTcbRz3V/W2s8Ap8dbsg0V1SE6KGVXUxk52nsb81K3FeqxeIEXBd7cqiNMKf86
C9OC7yDPBDDjD3BI2yar5OuELptyODE4Hw+7FAnw8aTZM6YlnMRt7WP4UUmVO03hfCeWNXl8v5xX
7OU+ipS7JEsbe/O4e2cyrVUziM+1mANzrqxBVcpt3aErKmSr1rD3qezRSm+dwQnj6WQwNP3Cf4bX
AGbeC4mvxkA2t4MUnEaQhbdxUVbJMXdRZqvAwZE2zljdbuJ2X8qdjkPzftkQS4SoWMfsXDN8D/CG
xp4myGjVlVoN79daRbQUKnKjIQbhfp81Sw9aVUb4kMo6vQFpAH2hcrd8Yj3kIlHi2/6Uk6BghGex
lo/QkHqODmYOWI6pLdwkyDhSLtxc4c+pcZQJTQUy8u7wqxinqZO9n+KZBu1ZKevLF2RpR/dnPB3N
UsnKge8lSWa3boq3wwxT6koAxFZYb10DI7ZQbAMA8e74/XflUUDFSlNgqgj4SX4DDkQfl1x/Pnwk
bHTZJhXH40fBCWm9NUogo22Gt9FnNkDjo3XdFy5SO9CFcbTYZ3pCBwcbvvMjyjIzIkX9kQY6BMNj
bpDQlnLhYOgEtC+Dfs0ejxkRLFpL2/oDJxoZJkozPy51kAmqb/CwuJ5ppmQfKihhDOR00NmEiaIr
CvJSqfl5u4zXjy7dWm8bybxlxds9VWxZRpVgk43gccWTSyIswnnMvU9/BhqylLhY6rMFNU2ehM+k
zIamowVMTIXrWkJObmSADWfRXyRZGkFJVIhX6oBeuvf+Wyl79TzcbAu6dLtbXrAChbxPAmKNyB7j
cV7OonBDd2W4YHELfBmsV2EnpLd3sxb79XwKKBXHL+8QwzX4rfNoLSQWCuXkLy2LznttskFdVTAF
SBBXS9R8yF1vlGMAFdhKpW5vTcTQatxhGVKONNo9W+BrFIrF1HTfQxDevIgGur6gQLO/uTErLLyw
W+ITghl3n5bWSYEbVmNJjSh0hzNwlE0gecnYrYWexlGWQsNIQ1riy5ZYmU1606dblnujWUql47Fr
i0ABJbBUCBUHh6rJG1eVkmp297zbckm2Yu1n5Y1gwNCgms8dTd2GRbGHmVq6/Bt1BA1ZtzPdd8Td
oPv0M1qpdgZbfJEGJrbGWjPC+e25qJfLmm3xBdRtIhn1q9aE4bbEaDmF8De1s8M9Thv06RcR+I1r
9Pk7SPKPcrtFJOBEYoLTgH++KAUrXSSxGQb+T5cvRsh0k00gsYYT8FloQAQqx4bdHFbyjLg4PbyD
yAfxs+tTr+GGSNoOEAKUPGHvrnyZHiWQIj3eqkoqMm+84nX7S+nA08n22u16AURB0/jwwZlpdfcJ
WWU6/Y5McAZ9Puozp7aaHVkzdXAmO9dh1CSk6U4oQkpI4vXzKZQ0qRS4BO0m4ck2SD8VYeRNQW4C
5qabpDujwS+ML/f3WPmh64JIpdNlmtve0YMRkXYyGKz0RqU2GbeBPzDPGfhd6oHdeiapHB2k6bL1
hFgH2vkU1kTtytW7eQF24+O52aQgy/+AJHWdt+6nBGgpG+4lxk1jnSdeESXuGknRUPkGCzoVi+NG
jyB7Wrh+eu8s+GStK50nyDl3vIJkEVN2/E9Pa4P5CV2Q9l66/bPhRtjQsevhdkSZHrYCSKlGHzSb
n/TBBvBkQ1ldEpcAXes1fiqQKhbU9NSGYwpFksG+sLZz1WtbBBFK38QbmrMkIsQ1v8Y5cFmoT2HD
X3T+z2vne+UW50LAWjD6bgMM03Q6X0V73Lq9EtEJxV5kf/1HMbWHXkYz3dlbwoJ48PxG7C+PFRNX
O5tWZzzjDpxfP/vWdHMJZ7osKKTyMPVBC38xJqMkKPvAVuMEfiVUa2TTIZVhbgkz+ugGOvKmneaV
hiK6iNNTMFYFFcwY+d8EiCmHw6A8UMyvKluBqhJ3Yw1wK6Coe43kbolao1BFmeH8YyCxmyAfN1Cr
VETDwqIhf1m/UoWrReUMGYPwtGhN+YMJuMJqhOBBz7g44zTFu9kqlPAxqS/2HeiuaCJ6RCq/hyra
2jnEJguRxwtm9qxzeANY6Cv8S/N5XCL7JIrLsKI9376KdH/CnuA/k1hF41ab1IA6j+M6mxsfffmu
ih01hBBQj12R9bBQnXoiL1fyURGr5To88iFaNx/l6vyzQHE6erv92yDciwgAxWb1mvRYyvIDLkYN
jsBlzrxc5BGuQ4I9VQp5Nym9fmPQUpzttGynCpPktW8uyamkmIomYteFtnYl85iNtE3lLZXmIjLc
9jxJg9I7RANrEdcw6OdR6lHuso1OYsLCVB1HHpiVeHwDE/JMsiAJIBHhhwoeBAj+02Z7Lvl8gnlC
GMOuwrGaKIUWWm5Re6QsoklrYKiBvSEadcqt/nFnULu+4SochE8G9VClus/V6e9mk0in2AYO+1RG
QhCZ9p8QzXBbbvc5NW8+cLiD0vZLNZ5vwHKKGjEGUl9vyqB+VUyZ2wZ8PoRn9NvHd2Fd3fmZHyPL
BlOPvEYSBM9g5oWbz+QE+T+DWmXrZ5FeoOquTSrJd64T0UNk01Mk8h6kGl8qHK2RRirI3p7e0F2B
ClFNShzJOcHzHYJo9mKhMYb0cHggZMwQO9euO6fO0jArreNG8+6g2Zn6y8HtXCprdA98cizMrCpL
IkabvYai6hP3DzGXyGPhVKd9qkSZEEcC+7tuNpGZ0ooiyv+10aGzGlztLEvV+DmhLCN9jG8U+/Cl
WtuBXlAw2FEqmaHwY48aQDPT+Wl/HyW3gHc7lbEqji1CdRpRXtxxSZfVGYvT9g+l1E324B6iBVGR
ytq9/LAhbD6yvbG5tAEMTrhqDpsK1hePDLeHBVvWiksAF/ZJtxzQxLjteqddq0Tv2TijW6umR9A4
v8src9jr3dfRRNsNJW3fZRbmf5Ic1ZgGR9AIi60iD8Z/7VgAIq4EF0zLmovXg2M0fBzvXUHxeMUY
lYkuOqEMU5QJ9gm+aTffcQZtvonaqulzpFbZVhdZwfTMgDAQpcq1C7Wok9yOnezpGFS4MDUNj5qq
xJni08K+FLX3ZE55/OIIfmLRPD/ri6egn1nmgCGmkxyp1o1InEo0Jfhoe+08PPWkJCDiSPszShWT
XbViyW0rTLoBiilxN+1wotn4mt9y9q4QLM6Lfy2wdxUI9hzCRyrZw2LOctGqMHT5WzCn1esviM4k
QimzE9jITJ0G66VZBnOAobchAWpvlck7xE5bNOLWM5aL8gygUjks6fNb2/Es4fidHuTdxtPBqIk3
HkEcbCSMTGW8UeV4zi1P8A6g2tfB2Zo6WF55RH/cbrbd/NALR1mbTH1Mi8ByyvWze2J0HetIoaPP
foU6lfpxQeRtDGMgLjC6S6WWHU8tR4YeJO+DHkuaf4KInmEiGUTv8fmJ6xUpmBBS/DmZXwlqvh50
rG+xJcSAPPkyNU9m3Hu5ljWlYAfm6zgWCwdK6HoUYVTgD+208dJpLPdhETg6oVI5u039CUAoDZ1u
e32a/cfdV89+kxzlb2JhkLl5DN7QRCa+8pUKY4vMZPRFclV+dlH6k0nA2aNIcKqD3qk1hSR5XqIl
Ovrmt5+G3szs1dTn9O4siT+hn0XkzX4mrm4OSuxppyGEoT28kiFlv6hjtdNHB1NN+yR4WkSlqK1O
+sJQeUg2+jdbYvuoIXswAQf/iyTlIiZQ0/OKsnVphFWC5NS91v0VPS6njGY2+P/4jlWmT4/Ox8aT
fg3HpUsKMugWUCdA9G/NV252L3KGrnNMhvDjuFybEcHdeQdVHyg2bDVoQdvKEqRisUl2X9j6NF9j
JF6PD/ShGw/X0t6IYhGXjBYdUDwfeRc9MXn4HPBIq8DQpjTaygGceupsmt0SbLy9mUMOCZj9TuL0
GY6LKi0ofwzJNfJpHVXfcECOAnky26D/s/1/y0Cu4jqHe6wkOtsmUnwCB8jU3lu0xl3t4ZaygdZW
FIQ2TYCQC+XmPFk/6VAE3JYUuuwE1HmLQIgGOL/vcgMcmiOTNyM0wA6xnpgzNsbxkmbULLoD1VG7
r0it9KgtqWS5YrDpHHgKTYBavIVxd+8YVsyyCKmMghQfXFyYP/yX8a1K6OwUZyLONTObWTV4O1k4
yCt1jfQnq8L6fmUHYqd/mJaoOYfsYxNdJ3BcjET9zbJ0umQkPEDlDRjBgAOJAAtezV5P7YwZ9v7o
YHKTpmCVb62tq90yQe8xvZXL36nJcZv4DsufcZ+yHr+MG8j2Q2BEAG5WpaewsaHCONNSNYuoG5QY
dF2K7ArNbCQaR6ISsvLTvYXCOdjtEw2EtywoTgwfck/TsgkKqOwDR2RNgCPpAOgjAqTYv2wf+mcI
agOf4DnkCcGtJP2uhsohDhv9ynRG6TW6gmwmTJbxpfB1fPBq5sq7DRTSRpOOfkCGLfm0TDZeYFVY
25/jWN0SKAfcUtb9o2bO7x0r2eFEXFkOsa/pni0c2JoRy6JTzZ3cwd+5r8oSPCNpj93moYFgDcy5
OYQ6N96YHWBZmaFSY5ZJkhJ98h7j4q7qU+xRPiZ39wDOluySfBucPvafj1aLsmIZO3pMg7IfoZEY
5YtpN7uFphKdR6NZG9riIrGIsni0K3zj4RY7rdoTpCoVPIOiHYyOXGXLOFGZyhLItKUSkoscLmfh
6qK1P6WGX5en+/OTb44U/9FA194g1IRUpQUmEE938e33YGixBBns2DzhrQnLrk5sqUm9a52P9u6j
F8NeDGgNRKqQ74byEWiNyz8OhbxCRHTma+0BJrWeBbcVKrE/a/P3dKNjAJa2/k1142DaA6tKunlv
kFNhJS9ZBrzaSIx4nMzXnTZBHZyouXfq5oeugcbpBK65JstDYzOXLl+WlGnfOmiI/IUnyC13OzK2
dfTAuP2FuIWnEcgUyoYOhgEEwmuJX5r6QKTvIqBHA+YKQy2+eRAt5MKcwDXy8GjrUtYQG5EZcedq
M6jJTOwnBZ7bwKMrW55WkuD5aYq+rpqXbi6Gq6o7bEEf6HPdzUgnvFf9L293+ljpWWev7sYF5LGW
PgyJHcxHfODu4FecP/vY3N0N49h/4hNC8hQeC2W6UVJH3WodWszb8zHFCkgQ91mleQhXQjKOdXXJ
DV6dERYJm2jNruUklWNQ9LBRqrlqQ2hA45y9RgTUlY7CdEpg6gPioFWue/g1CrG3rfXgJknJRrGu
rQ3Qw6bP/Lp5B+Rvae1yBXhTKMIuLaIG1mVSjqpp1Vof3u3yFsQ51sMk24A9bJsrn6Hm9PwYgKDr
dVc+wYenh/1a0ywn54mxBKrtMAt1EDgVpWm6jMYPYC7l26hq7TsjmhBJGuMls2pPKKKCJ03JAofP
l0JKiYHwW1A6352QM8mW7C7XtytPLOcoHlBfoaC1X+gq+2+ONl36KV00un7z4BON6OfwzcJOhKSg
wMBL61dAJNkKU+k5QVLcUVrJpDCmlnfx3pPRNBYD3JgCu5+vJqeTi30QgEABfJSm+JUwUJd4Rfh8
Rf9/Bl6F5W2pjnHlwW9FWxluMGmG6MELcyaiu+tSbts8nPr2FhFMdeq7D9e75FEecykoO6kwfceS
+okmYT6afazhfDs7m3N5F9mvuj6/uBkc00OlQbjhsf7q5xdtmf5Q42KhHVZ9gyyG/RurrlFq6iGy
JpsgN82PYFxQo9tNFzf6NkIZfsm8ChwT4j6HlJVcF5FLCDGCG3Jv+D2W7+pH/1+RX5Y68NVipEDV
huF8axgeCp78lIwZnHDCRYw0TavrE88YWClLl0l4HdhzVA7tRPxNhk9TLzFbs8BYptG9Wsj9JZvH
dOoqSeH66+hPdudXlijVsA72t2M1DOUSL99aci9n2LtFvkDdmtm2CLSVgbGRfiQrYxjH98tQPp5s
sKI3QZCsUn7R+XN+vHdTTspGWylmZ1UpwnlzNWuYyBJonCWYcaq+Vh7s/c4Ql/phitG1boiAvXpz
f3sTI0oUbRGWUjMp7PRwlUVJcg/SGxrxIiyw+cLqZkBAWv04/tuUmlslR9UjcWmXyWC4RYFOMhnL
qaBq0OpEW7iXYg/PMx+WFCEtREwWuMTd7yWw5Z9bWN3cfEvZ/D2hk5xuDLAMYqLVtg/IbgOMGfIT
Tl1Ucps62EjWMxn6LQrbWeR3MPm9R58DkimHfxPjzfGDMNLEFWgN00b6ifgQOOSlQH5dR68h65WH
OUJdwhmerHgevq12Wl15d7t3n9JUpfAza/J5TzmCwELy5VYFI2z5r5UgE4nqEMkyubiqUNkcrch4
wGGwUhsc1JyLo52ieBmhdFBOdME3ugjY52H86BEpfFQvknnmQVppTGXRzFAzUeU+lhTaZ9JwkoMN
kHobgG9CztW90EOeKdLtmD/kl8NrHVSRKpi+8fcLNTc7+VYfAsS1a8W05K2PfHZ/NvGaYjhs6EKl
Im++HsIXiGghwNQp+rF6gkg8jo7ORkhUKKBLuNi39NVJYMrQfYciLZ7GBaeGfEQssq4tNTgNmy0+
NC/yhZ3+ZTWKT4Gb60+oP4NwuKvJtUS6MGj5D4b5dZhHg41MwDU6BwB/fHWMHHFGygAsu/wMg/no
AVkhyqef800k7q2aVOTmR8U5oIRSrFs2R8n0NHoeWPXtwhEZcrkJ4K7wuxpOdnyg/tVIENQVr24e
08SmjfdqvF7I1I62wNV/+RdG4vFx5Rjj8nZfQhnv5v2ftBZfE+YI+QGQsE8suTrS8Bgb0yyCRYqU
fv4UGlXpUwiBb8l/1SbgdVKfnQD3JSfV82XmAaz7SCR/f4kVVz4Jnfjl/YvLsezTSTNi6o9wm7sH
uVt5TaS1wHEfrF0dVzEx850R6gCMFWEK01w8c3QLwuEP+ieTYffyKaWBUpVyC64gPGMb1B4+b5I9
/bzolx9/OdFnifkoBIAewyMHjWPEtkuU7KI6bj6RrDewIzcLiu6zMmKlh/tMrR2DmANy85BCSzqH
rryOkNPGihM1NufmErFWV+HlC1zk5wPBytQxSV+RPinEFWPw2++gqlzqn3bGKo8YPSN/Sc/d/hCA
pewv+3nIIXNbNafcmJVsEkNNejcYjJzTjzxr3/O+/VawiN/dN1UooM4QyJY3Jr4Y4SAD56/qpE5c
QLijcEvHehCCEsj/9KsFDnzQNNNLVjmA66JV/x6ZiPQP65VnNFMOWgBwpTQ56x6zxEOC9TCBgtMQ
WQWoL/zhzdcWYOsyCpHLI37S6zYR7Cboc47ju/iSImqE3Yud2CmKQMrW3sy1u9S8XOVXbc8NgfIS
6a9W/NwDTw4pCkXlF9QmY0G54l+/nW/9hMSih2hHTtW3G9bob4LaCKea5/TEdajsDUOK2dpfLTIS
RLhf25UUkgnOyu0FJWLctq71T2lek2uUpo7sOSkQTN2F9r8auUCBr5GMtrkSw9iXr7XHNL8Izzp2
FE3UzhyNDmxP518M28J9NmqgWUAC4bcIv8jtARd2tgLgn8zvOVTevRJD/S/UjZ2W2zmznwYF2eIe
belWHbh3xMtER1ef+ofvwztK0LAA4sxc3hi/y1PXWhntqVw8x+Do2xk4rvDfCHCQmqnoQz6fD2vD
mXtMyrXkVbPhNyCrf3d4flsWrH1XPkDErOhtxDhHeFgLOaV+hqht5Z6Vnen9umcjIxrUEjmz7Wpx
GYF/2IO9ySdREcuh4FsBtXqf3SZbDTJZTAWuuXe8zy47EyPPwVI+0vzU6BqUwwJgFWxZhDaWzcd7
9q2w5+CVpOylm8zNErzeAC+my5VlkxJ75DqpIdeCvl+jRcIWwBkCybDnIFQqFfilmjOreh2U/EXs
d7lSr7QhI1zwwvRCeIKwafeH7vz7VEmgefDKW9OzXIw4PKZ4Ry3/GsdAmJLDDljV5p+eoEpeRAzn
21YCwNNB+RQm9PC0edcWWXeTzms4G228cN83Ps/Hv5KHU0sLbGSUKgjwcxjdsZD9GEqH68hZt5Dl
ZPlxr0psNQkxM4NVKUXdFTGVplhKe6fCy4gadzC5wj3uexVYsq7WmffLzeIX1pyPCtSJBVLZynqu
J9UVTvBggSrxzgVa8cu/PGK3faGS6HPyr04oDhdiNGbE6KuOXJwFdts/zgPiSvQL8zKlxucpqT4g
eH7uSObeg0vOjFxg0n1J8njBdt3k2L0JOYmax/gvh0MOaD1YsvvlaNGo5ATMq5PPhbEfmSPETPvf
Xszjq6cpsqK8JsTnhcYB2jn1RLYlDJdtRUkvtuWMsmc7Inr6CaXU6Q0j4aLHaEo50TIGpqG84fy5
oMJerjcvwy6AnuKhQCm6RQT3oaTV9MgN09fEPHN+5raXOIuYGXB87Dsq0/AUTWGPakrvPuC8bbKm
OVXJC8JPrKfbj86gvWbsn64JdfPJsXaSrdukiwNdV7Nan0ITHdrxh4U0eJWgLAtHYOtOxQSUS77h
eR1Wcijuq/EGG5lWTWNFUlpdXOMhRM/vXTUbrp/OY4jTPIinS7Uy1b/xtSQpiK2jfKr3xg2bG9gW
VWgBhxL73glVamoHUVIZjZU3U9TV7+ylqa3MOULFnlPkYeTQzpvQSqUmH+Fz4N7nxz9jWyl4VE5W
t4PpSPcDWAABM9oP1GuOwvHJuiPVrOuk0ZBoHmRGb42LOChVQImUZyFR2kGCUveEL+aF9ey37MK9
dCy6LqEMk35pEvLihRa4+LiyipiNoIdPS+HAFMt6qT4Gfykig1iFE/yS8NHSI+z1CaMgidVq/3Mf
ZSzq3zBifJvVlosLR5J+HbHO1+NjORNCFHcj2IYLTq707QhQxx7jvQYyd1ohZsBUX4aWtRRW+hQF
+RSgt62w1mj87lmXjBdNlSbrpfwpD3D+49xIqbjUKZktqzOfzkqdqQym094Xtmq3kYPfm6bY2JAI
/igISvShLhCAxDOTiTUfteAnBVQjtZL+akEDTo7VJAaKZQy2e0dwOaKlEP7cA7OBfUJhPdksL7b+
+XYRcvJuyt6OSqzqgYm5ZH00KUJWbJLwzXJ1EBcNEem/rnp5HTpfN7mZ0HRdE4Ynotb1hJ7B7TFj
xApzGmrEtbpdymf52duSSkl5uSc65BlwrqBHfZfLwTA+58+FnlkG+cECf79giCt435O4c/STPqhQ
FBJ6VeVmBg2oIfaWU+BePGrW4hVWCJxsmM8iG92CrK5WINPy7ZZdANEsU7iDN203O6E3wINQ/H7c
dlk1VSha40SSc3vPvJngNJh+6jSv7KzL2LhotB5Rr79SGNVUy83qJek90QhLLC3R1jVCjh3XHVh6
1/iP2eUc3DfwsN78gUKRzo+0ncLWYmLp5/WC1JftEqvRdq2cDLCfWggPOd96DY7g4cyTsemgpbKL
0Xhh7eAIsn8oGKqNGHUNANu0PbzB6HNet/ruSjpT2B0UZky0Guhhe4WkNHV+xvUj+B+Phy77/XAa
NgmMPVxS4AbMwP+7t+aEaIClGPxAQb39Lt31LZemY+wDfhAZJmY6F2WyolxTlLk57ZW/KjEqp1xM
XdyMkvl2zlZeySsnMfZhhwcyFOImQ6lvrGQJ7an3B1W7wPNTCebqm7i+w3yYVWggd7NY7z3HYenb
F1fDCdbWb5OVcaYvMYRRuuCu/9aBYHMY7Jmd1pHh7JDVvJqQYjitewhTVJa/W1faeGnv/JqQTrGu
LDt6EDmWaONkAL+7XOG8gnJieRXM5YJPSX3HMd5grMLYvsMIBjcb6zs5EpfwoFVX40LHuWJdUOF0
R99IPH9S7Fx2uTRo07SGTB8MYL4oHjdEp6VR/DPNuyKs+VeJ6ss6SjuFbLMYUVKirj1cE24oZ6/0
URpZGVoO9x7Z8iXJiGcgKHAaXjpzzb4XQNHeubHWirVfg6f0OL+KbhHRJ8DsMao0rpi0BVHM2jJv
TjoY2s6TXWWID2PoHthBTxOxMoLIAA3Ieab6jJ2MLNNxzvO5h3EQ0s4EzEAPAxFW5B/dWcj9fHaV
BmTsqD2U86n4OU9m8zFaV/8lJLe2rpa+lyCxK5sBc99PQLikYNjew8xqyg0EAM1mgr8hGTAto+XI
3tfXT8Fi9RW3Az1/q2yBPC6zLg7NB1btyMkHFCoeAvLsy4pJEHsZX25yUzBhl6o0IFr3gJTGP7/s
Or4RxD8p4F+6Zhf7M8NzBk6pNKYxBIbn+XZkqa5MjphdJT+dY/XsnBrRmRbxyLPgzgDXmf/M08Dy
U9fk+6n4nk2c4HKBGSWJzsmd0OEuKG2xxemqj+3si8Y+8KlYWs8c7Md3g1fHxaSchdjxpIp2Z8ga
UvSDYyQKQX3FJI3DgwSsxFPKe/lJedo6KyeVruhL7o6zx3aDGuviAMWYAiEOzuGIMlzxS3Jjzln5
qwD+CS0Jyzu/6El384vKWVtBrK+sYV2pDf/ctdpMT5j+Xok3NsSLMo6QGQOWdN43/Wq7UnDNljmi
7kIDJaNWR/zK3Tk34JVelyNhDgJ8OpUTMZ4eE+i4WXbzM8HXdYZMAldTR2UsKFBYPy8yKaF/CjSt
BzfPq3Re6L4LRnJqWJPQG1sSRqMCT6Ze3GQQK9xC9DkVjHX1I/yNZXYqjrf/fi32XInSFOTxx82H
ZKwr5KAH3MR572eMx8hnOm1sOk34XneP6jQXjr95OvrO707o5UNyb3eAAeh/DRdDb3YOAw/wSOn5
7woJeKgVo/rpwKmm74eahrmxVJVxHROWH5yiECu8GXzycgfVT3xfsBKRcYv3lx6a8rf9RXvFvhim
nTXiLuNV2taZIJ9XMsxvVpzgrLJz1yykMrvULkYaNuGAni0CRSWMD3ENktDS2oEiP5U/aptYL/iC
haBl8BB762IexEPfDSipCHQ8iOw6oaAnmdE5RBiDmmoO1XHmyML+wjskypsnMNKdsadRcaLYlGQs
1z/FDs9YRF4F/p1aaf7SBphignUDwTCkZ/pAWW8XP3x4EtjLEIqptEuCe3LfTRWcMCkBPAWxIN8g
wwEtfJGa0gRtZVeNd8/MmjdRp1+MPQQetRScCJVT6dJLdoBos7l4eWijBEN6Jq3Jecjj6jw+hsTh
aZ/5DqOj0jtOApZ5/SyeZUI9mrz5a7odKAM5gJWtYTO3Df6a5/mByGeqoS100P7vNM2Lx62IxuXr
MGLRWhFqOp+mvpqJCDC0xFwvkhiG8lToXKhANqMt2GuCM6fd9iMmc/w+2VAyl5EKIs73P58yc/H2
u8+8Ek/DU8YCaF60N626Y+HrO2yL4undOdjo+4tIWqAeLjaqBqI6EigRDFiW7NgLw5To8Eh2esMb
3Pavw0XZdPi2wJRzNwNskvjnBGPVZMl/waGKPeBKFevKHiik2YMe70eoRYZuTM+ru6eyWfbn90Ha
WydjHg1h/mfbFOmRxrQQ6RhKjXPNa+Tzk+JdIqX/3+Zo8pISYOvbMebW3/Az8LOoZ7dcbhr+qEhk
4c9D/+PMQEvXs7qD3xIhHFEDvwE5aNeI99OMlzH6mjqLPiOgg3rqlrxIwfK1oMQF3i4QHJ3x+n9M
mxkC17e08EHtFUOiDE1K7HCU5LFHgAV9stnHVyWEchOBKzaYdlCMd2xq2dnAdHuKxFavKx0o3Fxi
dAmc/yxoUzybNA0NJsEU55iIq8hw2bWbDxUF/ClNlGkVWmDW5KpemapUKlXIVduP51y+ATuo41DW
FHsUQceT7mpJElmW2X3OW8ixw0bWhOgNDHDgClYymAzZUcxapww8o8r5lKYk3+TD8+2dhZ1pO4QB
I35DDlPiJdXpmLAHBndvMP2FsKaGnPgEeENTFEAfnaIETRf1KVz2TA6Mm366pitufBBJWiM+6p3P
AhlDEydRFA+eZ3u9DVBa1fvQGu3fmJ+wg8gD2HtuvFPeWy6giYQM5xmxAi/SDG/uz2RDXrx8WFCU
z2hW2Bnr2M6HQhBqBx5cpbqUIXSGwIabO6yH4erqP4JlaG6GA2UMZpEMjOebTLTiXQh0q4S+4v0u
sYaB+D0FEL7jkC6Gesy9uHrFb7fcmUc/f5pYbBVJ4rPn+qoeJzDHdgpJfKbz4gkm2XRfzy9ABAtX
oEXrFIUfdazXo4U+45JaYAGpqatI2oVeCAV1MR7YE7s7sJx2Zd5UlBV748lTJMIIfDw2Q2BXC8OE
XTbxVbKhAWOkX7wrofTMV5SwUVXP95+VCk+CFw4BJpuXPpM58HP1PZeeK3SsOwPcauvln3TfF+xq
HXn0+uXG/VqUde768o5xZ1/vSZ79MTWsw7thMg4DgoTSl1F4Cdl4G3X87pcckwxW8NdWrfHnsoZ4
73UEwC/I7FIgyF0r9nKcs/EJ8g4V8qy2bYeiUyapmlapDj6SKwCIh3i5NZutl3VqHTYa6PPQtswZ
fAv2QmnDeVj4Wc9HqDJW8xaADNpSkveKBGKE0l8Nv2ImTdppB0kPJVJ3xeRuiy7231+Zwpf11UPp
7kSGjQf2Gt44OzfzCYRdfM3Nwl2UtvOTDd4p7qzh4Z9IC3ewEaFS7hSRVYTBzhiAPHpcqzS4QQca
glDSfAdzE5hg+CxkTD8Y8gZ2PaFLRlHOTZaf1OZIsjr1drbM8E8xl1rrxF0f3d7QjoxCyZQg7Itu
3+LvVBnuQ0dOTtbBS6XO9sIlYdnUTZimo57QzeFc2vgqy1r8B8/nnedMl96I7E3bSO716uQ4kewB
FUAfrA9W0R7OmmJUq37mThlwLqZ8ZEOyUUwyiho0Pln68c3OcbhK7ND4jLKGpEZqAvp0S7//di8u
sgQFuiOuLNbIm6Qu9ytVr3iQotvtpe/w/qKApbOp6VCKI8cVIUaKloFrHDRQzRS1n5fCjgI1siLj
6Xv47uOBl1S9w1YZJgv271SPRKs2XxzpA34jlOUjiUER0SF2DDFt05m9o/Eu2BxgpH93DmqwjX5K
qgDKPGxI3XgxwMUMhyF0CbSu0IUDKFR8GhPIa7+QlOEjJM20zlHn9pAPaDzIb2w8BhsrHXBZEzXi
YhSnm1Gt4B0GwIlnMgprOOKDMuLaGqAkOUsYL/6eTAk5S+0zCRvbs7dgaHY7LG0IJXJgWx1PrMbc
e6hwKcbSiKCTOhl/FOJONhMvFBn1L6IUU6RqCTWNTuyxjImjqF2zjOkmevUJR/v3LcfahY1U8l6Z
t6rsSINOCaSdm1fcQTPTPfw5RTPzrjtcw2Z7NKeCCndk3B0NjLMScUoX7AEdNb6kH4mo0AT8qy+2
Y8+BV36OQbhfI9IdRpDxrALU3YV5he+WTwut2wNUtYRmP1tAatKVK3K4ij6r5AOOCRHAlXF2OW8l
E2V2I9cwl5T0LOe8nj0L0mQMjIpeA4MNhL1b81NpVVdj9QmYAGNk73AVG8dEwnn8OEhyHG5BF7OP
QAwOMgLYFUMGE/tNmvw/yEK08oBxAa3JX6SQqTwqH0VV5h5jvZ1GKEWK8ZdV7D+u2kFt3foyvBmQ
WlGYPVNFfMT7j2lRpQumKXr4VrwduznpNNmNp4ePTTpCTc9RK2U5kNhhHsxZrtffBL5iowZDSZ0A
h2SxtPOaDwtj+mUP6KgqN+u3l9SOc/BUbadi4qcXESChQ29Eh4XXDx0TT+l0cj+2mY7UBK1okZW9
VH7wpT913WTliLmlapv1s3HgXiGR+t85OT16NMpf8TinchVW/h2tKx+OycozWR/tSc8YhWeyoRba
KVlCJGsXZVaD82e+EY2kxNEfv9D/EQ8iSpxwIRSM2KLqasxsro2Cai9TDNANMyoANlyegKf9YHow
sluuIatsoNDvj2LJfdSe24QDA4LDa30SfSeXP2CJm1SwJUXu/EF0mrECCwKsPG8T74WZ0eXuoGhc
UZXFPndLXuesHC9wgIY7d8skLY51VM953dubBWEk6TL1SKv4Gzl0dZZdhtMmSmq4r4ihBzO1v5mP
brevlJ7Eno1X4GjYG/jfX+1clzumu/rTKknEiOjxrlmAjuQcaRZMtfmmtO/f5L9UM2oSMJu17c1x
E9TFOuxQzcsPonITjG5dfvf6klnfgR9m2F4GojDH91D4EKXlQSrCupEmdgT7hCghMTvBGCm1jTvQ
LX0hPJ+mVuIlZUhLiG2ryTfDtxHrQBYW6YYLdWegJT/h7xh+FNqzevLQ0ZJBk6QEgRReSJyIS+Hj
b/LBQVuh515QOaYylT1X4zPj1G3sG0Z9lOEwzrq336z5WOXLAZC7kCEuRQbZpWcaF89FGshCsvtL
IfPaP4jyV74qu6bWI2wkuJM9qmIfoGUC9i44gSrE0u6jSjBjdUWG3ueAEaEvUAXHISdwzaJ2VZnH
19otBMRtOjBG/zxvmaXn6gqnnvnKJNuki9Dska6BSMp47EALY7ru1Xp1jxMVVOsYOEpfgZzd+HyS
eLk3bKgefMNOqu+TOtC5B0wzq5orU+TprNykeGCcaCsFVePNAMBsFxXjmxIK5rOFMbuzcPMF6o2f
NajWFYoiYMfF+/5g8Rk3/D2i2rTaB8x0bDdCTkk35X0FBQPrbdJNcU4eKVBgt2Tqk4+ytkHBYWTP
3E6xeWtZXeGWcj79KT2BPuWQH1HbUtOSu9sX3xJmh16CW01fgsj8DuG413hrn9eMtk1LcfC+9eeM
pfMMrnrT0Cx2gTiGoD9HruiJRiGnyvwYPF7XUj/mrl9vris01SZekpAVUokNPspJgmOOfS1wjWZJ
rSuU/kdfR5l4INfdF9remIDh9lU7P7kWPia9HYhqIGyRtfc9eBQXJfeKuHx9Otmtzqb62uWUX+Cn
coxLQ7MrkRzigcVanqrQiC9y7EKos2zQ19QURhhZ5E9pjZ9Unlof7Ycry1uX49/1+Uiaioi3nFqY
ktw6PIXzok3ontscORzBjA74CVq2jj0n+IgXEf60rgO4O2wazGvxtvPYKY6wfMqNn6y5FL3hrjHH
WUtKVcJELmDCloMLeq+dJGOIsaEu9tOp7yAZXrNe69k/ni+lB4XEKd4/bhifO5UKZZzBNYlhkULW
1X019Eb8YZcC7PvxbLIzc+DiifVdk/9LdsENRxpQIKUB0Rbbp80DH6hjm3rJ74A9pqu1tYXFbO+Z
KIQoDG/NtMTodvfOFvq9EiCNHOfx6AuWvBCuTCdkI5IIXzauQshk0nPq+6fzjIU0NDflrJ8PUCWz
5+ZZh7e1G69SIUEgFTB5y3Rv2wXruoW3IaNwtUYI4AdWFt0odO360c4azKwgBfOKPllONSXc9Xjr
8rOk402MhQ5FLrnCssqhO3WLjg0UTikxoHV+yuUE4P36/8Zg44uy4hDcC03vNJddRtVQCRsr6l9V
SMjspBJm5Hd+ohPEb04qYnZQKqrRgwEJWTjm3m63P6pe5N4aiCUOt/ndnuHpQXkIZfYvuD5ez9MU
M5/tcVLG7RJP3SRiPPYQuS8Acthfrj51arJ1vMmpGIrDQGfmamMxMblQA1HRnU8VHgdCq24bK+sn
mS9tyba/uCrVAMN8cS15Q3cBe+EFsPIJlZo8lpaaFDCs5gAZq31VPQwRkGFUO3V1vW3T6MoPNLcM
OxyrlX6EV58+hbCtix+0T75VVyF9sjdxTx/p7U6kWKEYhY9whq6Ge4vbz/S8YlQsgC1m7ib9GGak
rdj2zXew3890Nnh4idDha1K55wW9aHmDXwQovA8QeuIhwPluoMdAk+shXwRjNHsO9KYMWWHfTsz6
LQHi9szrsCyWYPrN/Ek1UCLFKUOAcX9DCmBaUstFpKfR5jBw7RlvNxUXkX9CKimmGCKONVNiFiNe
e6ai5OG9IFahnd5CVmh488sBamXAFMJancjMgy0rp25Ydmhz2UfCMaqw5MagTbXZNVg1cu2WWuAo
fp8FTEtYpPKIv+ua01g6m+D9hhm7/KFCCRCgVDheFkIqV/H1hMqMHHhEcBIzaMb2VwozEfr16Ow+
kioF/RzyoPGW+GTC6y8Yznn+MtCltBbq8gxTP+etleUq+6hA91Qb/9ETGPq5OVCyVVjB9ucnAGfS
33WviSnw1iYYwKJyQuYZfiyOMciwaUUEgudev/vWx8K68GBjrI1kZIyVFK2CSt8uzyuQwY2nR4Rw
1+nQTsZVuZ2KLj1X8fKR9cjXO3mlP2v5eDggHiU/HORkaoHc3I16yHcKZoMYbY+X3mCIXl7e9ikF
luibn4m1aPdVR1ro40BlXFH35cuqZFPP3EkRVM8I70+rbeDF0HDeOLZJ+a81vskoKwJDQDR8yZU2
kHxFngrcwCjRo6g0rS9MzJWKuQpdzTBoeMU1x9v5LD0/XbUord4pM349gLBGdp2UzYsjbxR9r+0D
Q2OsY+ijtkY91HNEQgTxZAXErcM+Z8i7JxVDsAnrPY/NVSWTBuEZw2XXeIqcTiM32Z9jCTX7MND/
d3kJE5pf8helMWiNM9gMYbyKoWqUlwMZs2RMeYRn4+MMN1NYuqmksBYWuFRDb/nnSRYypFkVVWNe
sZoKVaqWEDmSeMt3eeZHKog12d3TqDe/IgJc9DySf+AxuIFVreqrKqYG/1nR7p4c3hMEI/iyHhxW
JiHZGuMsinc1OPv/sIth6IkamzRPW2+zobkYhCyLS8cK/kE8OnKjpYvKOVED1EvVcWx1x0JEJmJc
Cw04Irx9O7dp7QBF+Lgfp35fD80FpG5g2VGKjPV2jtdQjU7tH6/2jWalIvAGNaBU2339Cv5xfV9v
gU9yWitHEiRVTskXm7gO570qDa0MV7fYlugDHofvFq1UF9se0zzp896whuSzEeHzSeOXC0/uCnM2
LWox2ga+jKjv07qb8V+IRwKhPE1u0KRq3BTHFJJISiq7b3Og6n7Nw0mfI7y+luv8rcg4hk4daE7/
hZAnaUph0AVJZyyzrDYMU4wqHPNpyz5/lqYit8aVlHsSKT3V6LD6xItpxSt4EsH9rrayrSWOf0o+
8Z8oYn0JMYspWzo9kG162OLulYsflyRVnU09e0zIyboNF7A7e2hSR7pgPPnKfkoJyJEYYtL3yumR
vMOUM1kReE5EVzZjN7nMLxah8Luv2yfke0vZXkpKbN2sL/HHpIX6Yvdi+SrBzReHbH8fJe3bV1kU
3fC8GdvCA3vGEVaAN7Mw2vWe5Z8kFBw9V1wOa3cfO78ZNrvSYfyH+23HgA8ledqOKRQed2mMWDyp
rtjAsGbAspkmIrQoc8Ge4U0h68ExU1IKGwjfr2IuEBLMsPvkaLzgUeDgB7V/Sj0uyCWDXVgcGnKo
FtDtPBK849Mtik804GbH8cHE3204ZSfHuw9HO97NkslOzUMv8Ko3/Z2FfXY5i8tJo0BJqRR6UvGt
IQ3X65HsHucOuQGWsLLhNPEtsW8PbfkKG3JrMjh/Dw8ubLLtO7HOiNQVHi+SAKJ7JqwYGhIhm9Yh
8MeQ2HahgjH6pPVD7wc+TJLjNrEGbWVnvrb21JVd+gqi7BhcDhSGQ4fd8aKPp7aeqQcoQJth090b
MosNfZw58h+S6yhutFkAIxHK/nihlt+qjg8oe/zFUa8i97rPWsTUs3PqW3M+v+bE+a8sND2Ucy0X
CU5U/64DzuQPB5vkFVB5Cx88NlNB17VlQJvVVPWXunakcwAf9vIDLC9x/9bl6onbLA+mBMNiBzNX
EkGCJj0E9eRJL2jZBWqbmMOBwB4B4BY3ZzG8dZU8Z7UDlC7snHaNDpDCIILJW2N/671HD5oiOPhB
A0lCTHHc/4a/aZhTajk4w6c0rsv3o7BlQg03XYpVmWUoC3zun76m+QKKQfQvem/f0+Xcgdmh5z83
OcJ7GsFMkixfI8TZyuBCCxWe1N+uXxZa3J3wU5we6ArgJ8IVuwxR2fcmYZSFwy+XPJ1Dt1jovUHZ
m2QBXyPUGUGoxkIA1enWzNEd64/Q9UFVbcdKvUPzjlAcoBqzokbxuhtuxIXhIJyH+BkYZ58RRpyS
sKCO5bAGfOEhwjMqhFYfEp4pC/92ofePFVcIsOgIA+NRVeZFnTBmfUx83AQ3PHdopmd4Oqw2jfZc
NjwwLrIdcnFX+7QsRK+vap6AzLCyxulVT5Sc6utOZJgudamOahy07g8hbhEBmiPg7pyXsSjqsn0V
Ydur7oMR0KkD0o3UjOZEfAP15O3q3BSvvNMbs2wT+gWr81IIbAsLm58e66pAMqPsKxRW66WCneWE
Y2mErpUPLwHteuM88yRBOqb5lS+p3NiG/dJ5f6DAxNTg7wKulDa5ObApGjetwL21CEqz0TiuZYAy
2U+OhS9OiKf2lvCNeOgLQiuLsxFRDqjROL0oY7m01hQ8rgn16IQ7l7v+ivKpkPwc73pb/l/TuKsg
i4Xb+6/mm4qDxuocWMs30eMEOQt585b/W9XlhMvg0kdD2ltEa/e66DvrBNIICIvE+cVEm0mpBswo
on2eTmVp81Pr18wKmKmGlSGow3CirGnIdxEm450SvDXtVU44RvIA34FTk0wc3RQGyrcsTTjFDFsQ
3VAsuvjJhNi+1Gnl/ehpxR3X4LADI/e0aRRvzzw2e6CbZWu4NZBBJndy6cYmLaEMDFrVx8VzZRmS
tEf/jODHkCuIfA+D7b1jtdiE4wVLTpd+0hja8AhtipE5KCQcW64Z8DTZ/WbGdYfK62e2UeF5pNgk
pQ9dMLCRppUUpJz7b6TJg4rsOiSHjV4q05I2ExtykXi6q8kfpMrZKyTwmb9pvWoXQDGGUFnZG4qv
tc/eU0SR+wqGZHS0b9BkkY856I2oLX2nWcWLdKCK98UvS3orKss5xou0xKzhXUyQZJGeN7ddJ1Z+
Q/+4VmYT1L6GIcvCtdgghoGFwkHAqkWXYNpp8uk8aF6uTEenRc4Aiz8lo2mF3YyXPTItIUFECFLJ
DtPFhrYzfMrwB/483rYLTyg3ixcKYXlToo5n7m8esGvD1ESyPL/qE7HhVoz18J9smXr6E53pNxDw
W10EeNCnc81TivhoHJMx6EIaMoXFX1Mv/YDhoSTSSaE7Nx0wSCaTu1OXumDVxriVOgrFtPAuWmGl
3CTForc9Aj51Hlq9pFAGnhl667iTGZ57jEj0vluZMCI3ekFm3FhkrNvhXBnp077q7UGs2aqBAiNm
71ueQOhf6h5nm5uMaaxJ/04H1M+ToqzsCvWviNeQRRHaiVEPcGQJwhPZfajfpgZZXX/kAPxVXTB5
r5ZYsXeQw26ALHWc7RcRhcyEmuwLcvbVe4wTPWsSIeQ03CwIkyfHt/fpRslNGYawMAcpYRs7U+a7
bYieikn0y1bn90ecsqK+PoBJw5RPM+DqtgtS4FfJtpBkxrA6ohCb4hf7QDcYA0L3+/ZTTi4ld4oe
xakK+ODEZ/BQThaS8jb2USdEnZy2EM6mSY/xq9Nl9HNGLhGuYtNkbaMdZnY1khyFOS2N136iRnfR
pbG0wxB8Zp/zLpQ5yW0fHbs1Dq43wd9nT2Goo0LGnqO3IYQUDuWRSKYE5e3JqEMHgclec+6dkEU9
UHXqm3yAUf4YbHsm0UXv/Iy53pjDGZiX7ALQzyDyqpJpQh6qi5KwhpU+XGz2I8aMdojsCto9TVo1
kEWNwV2BQ6RUHD5pS8rsCDGxY3be1fAEEvmMon3M/leHWvGUXa3R/9gvzZbSoVN5Bvk+/w3BXPcl
3BIKI1babf4QxBGaAD6pwSxk174Ek2s8zLbxKZ8FQmqm4dbOWOwpoyNHBAM6w8Wb4Vm1sPnYJzxJ
jiPH8BImmwoEUbU/L0fc0GTZgzoUBeFDF907LTiO+uW7MW/pSu+mtCrI/rbpNkwedMig8DCcoOjx
wGvlAvcEOp6W1dFIXq0qPS94rMUAqhUpm+WnxJpF3/Cp3R7gDnN4d58PCCbz8C/ragrImhwQvr8s
nEtu7/ldpAQoBpvFTztxwhOO9W9p5fzfzZ8i+4o+x852KL4lnGXYrNOEiVW7UkO18KwCbGyRaOAc
1zdVZyIcz3NueOGu+qNs7cWiWrMr5Fp1ieqdmMFakRi7ytIr+Ii1vha/X8AxwocfmZ+d2vNK9C2b
ke/0pct+i//VEFt56EL5SR98mqsNH3R22durkmY7/uqZleEGVgH+Drm2eelGz84AK0KL1KcB1sci
x+xvf/quiMJUpjCHszDoPE/lMK2baAEceXwj2nBDmk7emDa1XK4aA1rkW5hwsWu75nREa7V23BLl
Q+BJrdHZmKfm+FUBtycG2xvcoxuG7FuiP95aWpPK1p/osE3s/4rHvp9f69Pi2AuP2Mdl0C+EqcZ+
q7muwgFbm4oNw0qoDrROM0lbOFMnfr0EZMXlgvseGGNNl136EyHOYUpVBogxH4shNvcUB8CmCtil
r4gRNfFH4WXc7afePkaCLdxpmFskYdujbk0XC1b9t3y2abcQKpgiLHsyeiL96lAbMOhJpOGvA49M
5HwT91YyZ99gfE1T40PeZZOt1z65l1CG6EWmfF3A2PmZFpCx8YV13b4u5ugOTAcBd3H4iFu6hfKG
/2dwrg07RUkdfdzwJOuUw6pWrtdX4B4kR1oYWtE36GrkjBV9yp5xtt9mS4BOPIid/PR3UirMbdtY
FHR4tjauvMZJlP8INVu7ZMwGKFScY0N9vOve9ri/OHuYNcqQ+B/az68LSuX9Cj8q2vhHhQrRHjlm
APAOb4db2yxFX8Bbe92jUxaa2N9YhqGVRu8nXIY761gR14qDeh7q6x6F0YM1+NhfgdBctHd2kx4O
02HKV56AqVSO2ooBtghIm0o8fvkNIk2MWNXXUZazje4mpV230D+F4t1NM4uCdKsCKFrqPTJkSbFX
02ymcV+sCmMO4NEAlBfk0DRI3xxAfhB7rqot8Sq+S2mhdNj4DZGQQz+kGLrd9mF78T3ipZPJ65wh
a+d2W8UpAc5MDeNCvEHoWVR7mg6zxMQt1CIbdMwp0Tly0egk2AOMRysAoGLnOVUmDL2PnaSV10+G
5TCtQKvP0D1kOtiuwTBgUcvkCgLXCNrHOYa8MEI82iD65+cfZPS5KOwfHr0x/XkiWy5SkmgBPBGn
d70b9zrmNTtTBAdKTrP5EtQr23GzA1phXV94nyXkbpoUx7Wvje9y1K/2ECLkNavvJgAUnLe5L+d2
48RRCP2sAEeFVOt7Dbueo0S0uAFZAK0SPpnLjA0SD3qCzz33gPRsWZxl+zVR8DF0/NG6CnUOwtz6
ZIOWMpWNzaaQmnUbLrk3YEGOVPsQaAdtWcltz7yYc6Rfc35T27QPkqQIygl/xJaeIV87ABPrUzNr
gl5V1v+enopM9SKYuV/9HvzVzDtyNf1Pu2px5z63W17Oz1ORNs8Vu9KsepkkEVYu24wWruhE4YJi
1mWllcUwsdGsE3RBjiBlFhHhrpA+JjJXAux6GGBRV/7eGOae16GQ6/fMr0LAs4AeV094xMOroLb5
s7YjYRCAJ5m3kyPQUNDHjktK9VHAwhnyXYYCbXXbTTOfOw4fz4RX+/oKe785htcIhT0GRqms/yI9
yVb8oIOpmqgMhCe9O11rxsoVHxE6TKGmdTC+M3XNruz8PzlQJYmVOKNeIaw+1+aoOX5wj2O6pO9K
aJQoT6sgaYWsb/aqe5m7pBI4MM25Wv0J8RhpxrpM9YDUNWrdouVvjgM/mpWDZXhqFdKQNYqrqxw5
Zi974srFisnP/vD6dUQ8s57U7MPyhZWiEXNgSdF3vi0CO+Cp4B/k0d5ePn4B/KgxYu7YIZCANpNI
zFEqcCKnNahGu+qR4peH5gxhRucfYWitgZnCt70MkYjBA0+oGpEUF6f5FQE/6J2fU86o65uQ9SkP
GMe8mNp2pQKQHwjQufZX/42XHx8/9tMSIaVhWfYNqd0c0SW9l8YB1JwMH6GfX1i71jui9EwvhX1Y
+g0OXyBZlLy+IKCcZSdo2ngjTrYadCAi1ZbdfgVAJ4/V523vNuEIVwTihwuzx+ARMDOdQGyJQI4D
Hg20U3lgd3aw/HTvlM/RZJ+Pw3wN6wymTpro8Vr+Cmv2ZU5MEJF7MU/bPl6rPeHApNDvvZMM/ywa
p5uIH9OTyY4OUrAMNfSbJ00eVk32r2F/itmdvGAF4wweRdMTwzm4mUo36KbtHfnQoz64u+Te/drj
w0jm0vyIsathr1j+z2NQJxKQPAZJ4u+nSGTTIyaZczsjz7v6GOhLRhVNiDxSRbTupdR9Pnvu8Ywo
gMLqjF7YpDrBODq4B/aaOQMJClV1OcOa9RpH1irxm2Y8YfC4u2cu97PvV4f/8l+Z22RemJ/WtNyr
6i72e7AbCptXZBtBCkSIgEI7a7x7RtrCyfsdDpXT5AH/xDrKJ8mKkaHBTp59fxld4/wXkpbzTRsi
pr2J3cAisSvXo3xDapFIJqrbMOOpPL5BFnGo8MN+siQv4stfontMvoExmMe+tPi5bQIXMWS3XiAJ
+2+erZEdBIkA8fc50X6Gpe7kE4tkPF0Ah6PpU4XnK8oRjG50htSJ7M4FShycW0b5XFp8rgVAyubK
8JkQlCooLAlDU5sPRg+5q+egdE3BR42VJf0uY9eDM+cJKr8XGnkSSTUY4zN6zoPg7o31Coob8WOC
iaEjdo+12lvpgwv+UJRXaKnxFyafG6l9FEo6I6CKQJ0s3kkSvIyUJKy+kQdQ9JMk2JQh/894c4Ay
+0F+47VYxFy8JxGVJesRWV4zzYJpdXF3pNp4iwypc6hUTcVlmSpCvDpzpDHdqmQ2GCzeR9uIcEUH
9DxFX9W9jDsYa/g46ZWve4SNMgHeVRCd9OUPLUQHFq96cbDiT/hA02jJa4y3necVjF97xyZ4kPfP
GQGip3ZhJXLfJmBJyyickJSjwGxa4+nLD75ADeZlKJrQr5agWXghTJskR9uDN0WJfW4jJHfR4Du2
v8Er0j6sDhStNSugGpSFMIThLNGXxzSGm/aDKs9iWkH/q11Uiusw1rIDarwFWAPOtdQ73xJ9v9rz
ryskr/ySal5iei7pm3/f7t9OywgEGyGRatLqsFLGocqkRabwZZceKq0DnVnJfBa/X+9ygsbrEvit
7QyuplyWezlJsjpS+EhpwemtgqfD3DMzW4GeZfq5XiLJajtCj6eRmYQfLXjA+ROvoJsQuwLuqie4
uXpubRNmTbtVwvhqMXvoBv2tctxlGHREf4lnEOYDYAmSKqZ7xysZjpDNLvSFX18cvidh8sCh4NT4
qPEhGn5d26H4CQ6PL8UWpOrz91T5Pie6gGuI1C2iv06c/eDo12I1Iitcn2NlwOWaehcaaCz1XKky
fywWZs0yPSOwyCLHsFbkG9+ZBwctGDpfufky8lRQXWY13XYawcrxuTOAldB45GFyIAm7YCTwA/j5
86RxiDGuUV+fYLf2QESQ5ncF5uoj0HMplm9NchChWKgA/QG7uVfr5BNTq4pCXds0Y4xpkVM6IFTs
pRogqdGiTky9guF+l9N6A5VN43C0eyBEABTBEfvACYvcPuvm0Mkp/KgkVVWsDAH776hVOjU4GnhA
9z3PlourybHidL/n5ZpiLaW/LfPvLPtPobOIrmDjoSX2iNaDjigre8ZeJ5kabGKH1XUT4BpK1hRZ
nbSwvdMfAR3H9vTFDggj2Xvhm7rlNLPGdlkod5NsPOP4h6m7Uw1Z40oRkGDoFSSM4RkMnOy48ppi
vD3+tBZqp7tAV8GQSqflN9N2JAz5N6jRRlO8ody8PcIrawXDBXrOP5PS3iHo+YSaHKr09RbXr9kY
peMW/OvZ/MmMgGVHr3TviYYHf34kDtL6awP/j5eQ6VfGMCAjlNSoLf4mENYQOcQ4dhW2WRYEf52Z
8ZSchX54tFJNogq+9eAnH7+LCekiNh/UBzSK/Fg5d99ScGr+kSCOIBp1jpz+3uCuy88kdxED5zPu
6rq9vzvY6HQExNzHKZ2XB4QTHjparimu7QW775B34nnjpzCKXGlgWs5ADL7VsShCWolLRRYeKXhQ
n9AMxprbspTImPwsgNyqa/Gou8t+alkBA7a3S8xY6ed+wDkKla4jPVuCRgvO508zfcUu0ViiTVad
OfLt1tEz8xWPwIXq7wkLSUCYFzLQq5sTqyWayUx+oA1Ks76K9yfjMCyJQ/rl2vFOsEL/Nsxq7X/Y
fN5z/A1NnS6gho4NloOUMYm0zkPlMOgXqRk8jtBwqb98TWthetbGpV73TOq+TtfzLJ4tFcy7TNCU
zX8EaoU+zo0pDNuhsVxMKrvVZ2GyGZc3Ityz2qEwJXnjvQx21EMyrRQrm3qDveiyWsKbt0PIG1WQ
GTGU/EreIwnJ8Ps9leJnl6t6Mg//MKMcpEvAZFQGXWC/g+0dPuvVG15rFnCKsmuBjU+H0n5PzZB7
qL1p+XYRg69s50+rKwfC74yxX+AOUjfRuBA35ifG/iTACFKx7XwWasgWyOVx2HCCBsVgr6ASfHKB
plq7jiJMQwvPoTw9XPkHpSkcv79hm9+hLjeH+pTQhGJkmpHzpscJfUw81twqqHrfN9ZlkT/oGwcg
hz6L1UJotGtyHSa8mD27lj/gAfqTuMKmGZwOGYjaApYvm+CVh3z/Rbgf3XHA1CKOxvZnxSKXoRbm
hvioao06xfn3fAZXoZbD/bAEafO+C7otZVWPyYFssD/Yb4+YYYmWSpn8ko2BHLFjtFGl+E4zlgkY
rZ2JZI/818xML4RrcbE7aaNxtmaB3EEt3X+BKXlcQmFcCak9qI6rs0U+vx3bREa5ddv+zcwPezqK
aMTTS96zatO3olw4HaJr0fUAWw+rzBOsLlsFHw+Nh0D8aFVXdFuD1j1yxals45Sa+pxzGm3nKqP3
K/Dg1hGw0SSGH5gAOExWODT0jKsNjgkux2iiGDy14mTGhZVF3EQ6uTQTtuNHIzVXQ9kxSAje49a+
KNPGPd2pgynO9f1fco5QuIEyjaozXtlDAjRjlcbWZBzNgrlye7Z7ROw9cp6cJ+SbCiTXBtpXiJVT
ZkvvxPg3e7Gjrwr9TYkqor3GElpPt+xgjbO6AJYyRRp/l2VgQ+YPgY0087qj4JUzW40v6862mJnN
p82B99AjB6IEDl4bIUJMQD7w6ynLd8siHWoygkT36zlA5XmrgxKc2le69o4eu8yqtCQYarImQBAm
Loew8Ell5k6HRLk1cezBb+jNiT5N3b10nuo7CR8MAHNSBq1Ejdf+ahV9w8wgq14Xx6KED2do2TVr
kVg4bqmZNaTlLLGSXnCnYuN2dK30SoRDAodNtehXpXXaE/adLunplcjorDlcc6KbGbS4Rbs39lBm
zbzj1HTPyeLE6F24gMgAnD3pvlwyTUTNJFRrBfqBGUI4zLaEnhp6WpzeLk2tcoPkb3nLavdngNfn
ZLa+VWaMBOzSq9Em3p7ir2Nvk1Ad8x82XcxwINuWbRxeP66132QvfYLQ+Rrr5IJ73Uk8iCgJ1a4m
0wiuthLUg/J5zPjPO5UA6hUfHTa7mq836fEdwOPLnsb/A99bkvX95ZlJ4uBalF6OLVsn9LCWOdMJ
d35DiRDZboNTQu/4pMlQYU0MyhIwF+WcINTzLgjQwTGEnCVL84v1U/wlJduVIKj0ynIuZSAhOfvw
bjFWu56iCyCNhCmTXEXRPm56mTOFSgTxm42fJxsrBfMpkORom34q+VN4T7SnJutvUhzHitDr7Ahg
dksMYlK+/Ms+3ZpfQA6rgzVw9MlTD98pg5WaCMmBnvK7zNznIgezqToFfOQTA9dc+3BMaymmnAU3
iKP03qOfGvaprMv/ukoKKimZ/UOvsLV4RzCsJt7P4kbOYgBJxl5GixSGcBxyAOqujL/ru90RnWQN
cRMBqOTmmlMk7U/VO4N/CvSW1p+crIbsQglh6pMuKV7MB9Ic5xeO/m3yZHAc9cRKO8aTzmyGuSdV
vEgD+dVnPik4iwUGgPv+3x6ZdGEAi7f0w+5/qctgEK1s4kImF1hlAfvsYliYTpn0tyRK17UXLXvF
r47XCY/xXJfXB1+HskCxkD/8U7SHSRz3WmPvtETctKoMOQYIDGse/+wnk8DO0DTLX4g09Bgt93xs
QieKsPmn4ZkRBHnFDlFwQdZf26g5DPA3tkBUZUUTaYZUi7hjwS1mT1+FLcEKVlbpktUlWGgt6K1z
HsqOb3uUm9vy3oek/0ydZdXF8CBprhMJXKeSMISFVuAyVXcBgxMGcV1gjZHcIZZL7e94dls+GiWY
SiZRYDG1xsrNTJYFGtcFMnGfKV7Hm2kjARs5nBJHr1RsEmi4NxfJeH+rLJXuK/1gIShefYDfF5tu
HbTVM/EsbwcJ+H7vVE6Ii3dOKxLRy1f3bVMlJd29X2Lh8r2oSh0lPqYHmVZL+RMMmRgoimft3c8S
oM9yigovsEalkYf//ey5qIqgjAyXIhXCGB5MIi+DuY0hYoxw9vtGClHC55VWIN9flyPw04YvxuaX
VXeOq9NyAD7f83vydbjPLTKRBmwdPJ6FU63PMd6EEtjmi4rqkthAa43MdUzxfShFnMS0l+CR2gnD
mw2G7WcyWB2ZYwOprWG8qKZ74zRtCMN7cyUUwmt32cLwkGgzlIAcT3LzUc39vCu31l9pbsap2L4E
EfktlJpatlhgXsY/8hCjp/OHB7Kd+PXWkITzTKbPMrIZbPqWSpwKUR7jY67p7wB0FSx30vEY2jGp
uNRJYZpp/apwI59AE0bivdprweb3Y116kAaqrCZyOrPkrNPExia9Exqu0egaRqafMtmvJ7kFjUaH
Pjf1sq7tf5I6t6obqDNbBDM735tMLOo0tBDXvPsbcLOy+gBQLzLAG/RbuBZSnjr3K7BphfkY6Es1
2iMpWbd3vhJiy/257muRp6GCzZVEHRJNKm7WOb3HPfqx9ogMk5ZTw67wyTkQAAWY7PQ8vDwfLUT8
pARPj0r8pAadY0l5Ql3k2PTzcvHsSoPkBAAJ1U5zESWySgnc+zLPYRyOIPpmcWdl9WRJIN7sOp/H
gZGMbRl+Jiv5LZHKykQUXRrKVRFdj7J1tMIspRUVsJmuf1t5E5/aJ4mPpvEnt+CzqO0AIXhJViZT
wZY94S9GYPyLyl66Ylp4gZYBfd6oJtbBwfBrkPhvYOc3DVo4zE8Jw6dNtDcAd7P92oKJYSlqAGHl
fdUDWrGbPKLrw7F7NviYL80+pSQPH2ZpmS3B7F+tbtcloh+qySJHpORH7rBjP/0LSBylCI2uLeHC
tQS6EIS8x6md31fEj0e3GTTHMqYG60C+A7CGEEXwV3/3/e7I6IZlroQXlme8UBrxbJeVfsODvzWC
mLfDbBwpQ2jyvXPtziCUhdU3hoc6J3rLdnYnltaXiiZqaoFOOwTRXBGa0ncshyztiYkvRK5iSCEO
Ijmu+pb+Xv8+uD/eTfwEgIy1YikP7wpi9HDBguVeqQYB0dCDqkh83Pq+9c/46wkhNcMxE5wxCnng
9nc2HQrLLw2VhQbTR1gzWwl7ftp8JCo3UgINLa4KObfXbyCtt9xSqq0wjkpHgmZfvtzdDzZpwkLb
6a1/zzHBe4QamkhbpiaAKpqlYK42500TBvhTB8GncPKkKKj568IWRy2gOwhp5Ne3YRFZNH+1DbiH
B1N1MKQiTYdJYs6pvNCEpAMeg/5X4crBzRrC73hc83fo/GkR6mn9nKa3e9DcRVoI7t1kLMcYC6fZ
RKbbzNiD9OW5uomzohuQ4Q3RaE8kgyY5afou4HXaX4L+ltPKqxkAQfRVz/pZQ3XmMWYBydqqiYUR
Kx3vG02m5EvPp5sxsJat8VFkovdDFhiQ7LNPGeFax/gEnQplrznJIsoo4fAiwgQs+JHHENcfC5k/
Gb5IpxwXadB4+XkJiomd0wEIE1XxRvYPAo1ke0FfhY3lTqBSAU4rXXbvXVDlL4PcnxjBpdZZNdGf
BgEPBonOSrk5Axf7RUXtKOJXwjo+5KBIKAYbiDsqGzSGJ/H6hvEv9GPYxcKxxPvGci+z1IPVhdK3
Cp7FIydS70SG/Q0Rzhsab6oTiQrkPvJYG5gREq5dkx//ovyV7hPzJoHVKYLhXhyebeAoHuo0zdEi
pjrLcfnO32pkEuu5kfkNcGT6KYq5zX88R6DbRWdWhYWWP8UwqJhUki0FIrlioURNQNe/al9I2PWe
ui6tpJafCALd7r5tDEoelgB0B2PRui/usakDub1KBvk8RTaTQ5L459Eu7U/VBYCeVtEszXg3ZJhi
tUbK8kCtswG6FRnIl2dlnuqHxzh0wxIJvnTlrkVANpUYsbcLQKJeexodiDCNv9hUDWNDe0GRn4Yz
tVag0DnLn19pv05HcuIVA2l5/xK+pRVmctrxIPFPF6w9Nit5yIfkj81aR/Py7wbyKUyZBzEeU5IJ
zL54jF0HePyjNfuFyzE0NruehsbQ49OG9W6V05mUwAyxb1MlM43du/vzvTmeDOCy3FkdZBdyIjjK
H6ON9B5WhuaAsoBSnZl0mCxwzDprnKgmglxMqmSP1YqIZXsgno/t9zfUKVpo+sVsBpPDE7FbQoBX
gRbhZ1fFWdV4QxGgsAd+T0i2uMtSM4bDsLpB6nm/GD3rcvxAJtiRKUim6lUXZcnfCeSTYUnjxkm1
ysVrG1Jq71CLYKAgLCKsf5I1RoExQ33rR+3IbdiEjdCcRxLxmMY68s2NWyudSAw8fYjP7FS5YmUQ
aybla0h3sPIzpLRI/Y6v26cVqAildSVNCg8IGjCeZVkIFI8JVMtXJJrbdnA9Db4jr0zW1Q3nUBoV
CupmMozhTzu6FOHg8RNdUqlGqPajo5unGwsWQLRLZB8F9vVbUjlU3fsX5oBukkHQ1HbDwby28hf2
l08+QXXZQ/rX/d58P/VhSF7calZY8G0VNuaaAOm5TAIJ92SW4Z+1AR0kRKqWi7q2hMK88z4nhL9C
U1DIOnQvT0+DmKasaxItV8Lp3EIeFktHzUdLr90C2TudLICQdcM0cWaoDk+XLc8wQQaVnQg9hUjF
s++OYrhT1cHHx3H/shLoLEXXz27qJu+DC150fTbvlqOf+9ybP2DeO4t/EWTpWQPqX8zug2D5n2J7
+/+Bal37UlvnoOIvS4FjkXK2NZUC1recgDpdA68JMtc9R19I2zVE+HZ+UarRW4p6a4AJyn/1t073
m3gZpFC373huMZu8Yh+qrHrT+GFffSuol+DB1vRN3Dp9z+OHnVyA4mZXG2AqHa1knw6DCTHDzMqP
um2mf/tZjDUCPbQpQ9vv12ZAl31J8mSJ3U6RKleDn0fXkG3ej0ErgKEUrxfwptBrhNYHcXjLSn30
4mOyO6Qb4wjuziwge+p6gpgej8F6da0b+3IZUZ3f/SSOpmDUpWK/Fmpja3QFTY7eHnHkAfLsd9R1
827yq41DHDoCrczQ8LZiZKPYnNbq+WzxX6Imj3eCUqVj2GPSPK7VrzrqjdyqpvoyNbR+s3/OqvDE
FbFRgn/VauyWjynN4yFLafeVccG0FirKvpvQpj7dJ/B7Nk/PCvA9CM4T7EUYeNgflbgnRDLJd5YZ
HJxzCQQyP6JfmqbErpZiRD1TuSIsbqnRwpl0Ss/JbZqKopHbW7tkefztzDqcdDdze4AZxXcXgf8h
SLWpybUxu3uzG1atkFTld0NwW2qdf1vR5PXUibpAJK3RQFXOpYMhwiOHuzlvQyQMhkq56ENV36IM
3DdiVIXAoEgKCGt5nbAx5xzwEzwhHvoyhtpIWyB1Td5j9A+vbJceB8b8M2XiYUxkVO4G0vTcmwe/
VgBiM1Mr5osIIsr58BIvhR+hzhJyjP5/P68ToyYOL89baMHS7O3S6VSANbsrO0xmNrY8a3TlS3sl
6ztFeRO2Rp6oOlKz+OX5iKiSzdBBukx9/bfGIdA0J25Cs5HwFMgM5O9iwTIQilfA9DJQObGXG0rb
oWOFIiQY3VVVtw8aWxgCERp4jnVjQBYzARbBknUXVm+8AEXqoPBmUwHXnG6TkC8rnAjKS3nhgOnR
ZnbndkAqnD78SwUx+iC7rYvblwCr4eeLoFJ6SvatnfYlxK0BO1J/Xmk+apVsJcwWTDI14IkUqZ2m
I8NI3Jf/jH9yqZkXWk4qr7SjoHnuit/Dhl8vaFu6/BYNYWtZVnqlENPu1RZ5M4GfcR2ABsRQFUJV
hiQ2uXa0N1Sk7cndhiRn1wed6yilKQAk11cREM4nk1+LT7XgDPj8DpSlKKqcNb7krE2kDoE4N40t
7Dql39BAg3IOlesSdK1iLrehWzq2p0E0DYBqqTiXnUftrUe9OePphLkdRYjCADkypFtuf++Lb+Sy
OW3UyI/F1q7sU6toauhZXk287KQRc8aEPvuBuRsjVxlGbyOiweCKlARuezHx/xVG8LwqH5/bmVKr
25KijChmEQbxYPxddtbspjIYs+uhlzldFZUauBlv7Wi+R/E441hPkub3hi+HDHHDZXQqff395UeR
BiMnZBrnYswc5WW6gp8IvQae7Ycm43PJUGhbKbxN7wyGqvR+wb3DhLmXq81Ne5veGr2CBornxLDS
iVihZ8j1OexORiBJnmU/zH7WV3FSq934GTw7excvYTQjbT4Pcwf2gKnSn60F67fc2A1G7RLx28IB
LZcKSmWIlobDplNYcKXgvdEJ+kCgzpvPCENZduJgixkNKpHEvLRbdZntj2gsZtccjicEG5/VAbMt
E3CPS/RwCs7a0zOon6/DpryqVAtVOdgOqi4D0R79dt2Qh0FbG20LHYx78Sc03C0vCaFxrgAnK/gz
a5foCT9s2XQe+zEXSavu8Ptr4yalEGbbU3qg96RHrKBmrSBHlIRPRB+fBBy8ERuidpW61ZvD0I7v
4pQnpiLqdYpStkN30eAPMbYrwcRdN7THpL5ZiY2LcFWwh+rwSg5DRh20zVFbV0GTUWm9wqTjUvUv
CNg7ADbvY/UXe2Xo6jK/BVi5DFqKduVh9lhXqMxgU4unrV8W1qM+VnpqhB5eniDKho6yRmYgSsTY
I1yLuaNOKqahGCi8YJuCjF59yXCA5cPgmyHrZO82kmEeH6YLiGHuNlQQtxDLh5/p7xqjl/I/82RA
eJUBeoE+PeWxcx3NohuBO7TiiqWCf9X7qtp0H5+neA4Lq2QXzHnCwf20EeyxkLigkjST9DTgtspK
caUHVzJek8LcIcgKTb9dCH/r37oE/bNrRbQRO+V260Bf9+9jINJ0v218zJV4gLMKp5ZqrHMNJLQ4
xZUFwv4BSt/rrHjFInjMQgtKwHKMaMj9hsOVVXgzch3ZyTIoFAh99/+3HmAU6NUEjyGgeWAsO8Dh
Cmp7ANVjHdBA5oCqKsyg1uiLrEcAda3oi1P+PK0H5IagGQnhF2GIPF9bTfzAen2ugYXa2pRhADUn
ShAbQnkvr9UiOz52h9sgMBWuxPDjoTm5DEpNx+wl89awcwgYoPUoTiM5iFsiyQfrgKhrm2uICDNl
0UBZF9T+9Rw551A9JcPktqQJFg/4RNRTtigAgrnTV9j1GKXl/XB+XxdOGcZ8N3ElkO/QGFCoO2Rz
llACx6uzwUIR6ztfxM1hhixfInVuUoVdev7NoPxqtyZzPqqug3+gr1oWKLWxYc/GX0+DHYBLEiwJ
Ac8/TNNKtSmW3981cU/iL0NM24eJHEXw9EnDf7iYELGvIWGhp+C6LSJ9fDXUkgy4328DP/qUCbjK
pk9HFvAS/LQB48PplZmERU9etRe/RWjQeqVpk4qYSpuqppbxtdekeqva/TSOJ83t1Xo7Z8Y/ytt4
gOOEciioDHBHgkMv7MRZ/8IPv9quokaOpBL/T4NN1xFns5nNBkrfH4yIHoHSVYHLwCe/4x5T3ahh
7FY/fkcktgAlTMmcd5BSSzWnanTpOzHaZbcWrIlMiQSQ7LVU2elXc7wv7oBoDy+IxUUSdeh3SZgz
4s/gwo/VRqc0uEdoG7NHrVm/z3okfTnGpXdxpNP3YulGMtDTmhJw6cb1pJjmWdOWp5OuVj+e35QU
XzTDsNzR2F5T08Pn7xcxwOSBwwPt0AP8KhNMLQkI8erayv1plVj7/MKHMp0YB/Yo+v2MLPFmNyax
794wx0FSpRkDVYFTmIg1RYD/N4rfpu5dPlN8qC4lMmuv+AhrB7EQDcypFibzgQy9wyIXT/AN4hzo
zqoNG5eFzIw5hJt075VJI+JPRFHYgnM+iK3ekKorKtPPnNo7VHu/1wF4dURgtlwCQ+MTiUyelaZQ
yNZD3BU5jAPBkJI1MrSUPAtLEbXlEkNqiF+iLKX68A/+qLQh4Ggav/ZYBgmPOK+6WJ5kSdQbW+UE
v6dyJ+3BH7KluGrn/vCXAZiLdLdmLm2GaWeGU4X3cLCMVQ/pZgjoMHEc3Okl+k6uWRzRU1my8xcq
AaqIj08N2w2vIfhTHHLqOysQA0e2FLq53IA6URUgneUzz3k64uz8+l3l8t/NxRq+gwjly6Kw0oYR
Ll4QgOllBjG/3bkWbkl3hmVhcym47akNFaxEN7SLpIvcPLv+E4VsNeUJVsF2y+84r6V87qhHwiau
d4/DpafsOjdqvbpt0bDg0Vh0AhSQRwBkh7CjtGzhvVPAauozGq47UwnyqjPRnX1e2kt9maBX5gWv
f7TREcqYAASk6V2hvKx811Us7hF1iBktk2HJjZMgiXmC05044wYxQyd1xyurbwJ7u97jRlWmPhuh
3c3T0pDUJqtw0vSMQIfRqXtSyFXKYtRw8BWCbGVKvXKx6ML8u7altZokMbHuyimh6cPFdiWiKbAv
+cZjlCCkHDAZ9XyF3kXRpaCZjSeJglDB+VLmIbnIH7vo8ZJpSrvFnLGUTKQ9WCu2RPqa7mCP9dgX
+r3HueIphqT7E7blfiALsqkJ1pJaJt4NmnezlVUwOreYTjgN3dbiWmoseuwcHo1f+vBxB1WZnnq1
MjHr+sphC9SYNi6ed11oxj1zrexj1hfXNXh5M6Ww91Fym9+eSLNEp/MDJBwDN5l5+JSet3416a+c
K7VDaOBMDxyhJ8m9bkIDd+0tcfF3w8m53KYgNoG1Srf9TM1agDqPlRjwR86wpS86FOXsVowvkSOD
hxlMOo3VS9ndRGijvhZYGgn4ondx+VX2dNoNOu8ayAyPGT0HHeHrcO8ayHf8X8Z52kgpDAIqPNSI
BWI4/hZROPLv0xAUAKn2Nqi4Tm9spFPmsVEwUq0ZCUs8nDsGUbDzDYTpb2ZuvMhq1mQYpNWWsoOL
l+97ynUbCN2gpBLuNByJRHjcBEtr4RxDBhZ3AnxaP+DTenOdV2H5iPEuyLusbzZAivfWsCE6pRIj
WHc4GCXatBRguVgKr0vIpBzAFlWFKd0to/B19YsgAg9XKIN0jcKBrpoFum0DGekX5AxSvhViXLch
ljQgMMExaFPksKDpHPN5dSiPh97iy9mNxtBdvtT6/LsQpYNCBFYBC1rAFVInSdRpWfd0sQKGXNNi
CS2M0oVEjl8H5WcfgVIANZLl4qKzgLbXx5yHd2JfObuaKPFVLJ9RFJrn7uZrVCnKKyDjLm/uvInf
HUd3cAil8E2ZQdHQbLolGKJDJZpLdtyQS4BM8TRgOrlhnXetyWrtuiQeKpOaP+S4LjL/DM1HAVV1
lc+g4nZn/ul4VMPazLzDLMRPJuV5U1jAUglhsEyhnZ0SkARKFgsWZPsXYI3t///7R4w3wTmLidmL
zkRW6u5j3q/1t6nCWu/2ldAFZoo9rJC/9A6v9z6ZbNBx9ldyiKE9FnRayeTnmr0vDPKkPLIsowWS
zkgY2NIgj0IOeczASDZ/Fc6sKgu5upTaRsAlgixmcP0z8X52DAN1uAR5FT8bfzdOZBYBxsv+j8xo
2ApaRsBY/RNOVRDPOmCfPyy/doXQHu099nvqiAFQH7y7ucoDCpP31oGeCnzOeITUDEVRO7o7N7L8
eZXJI8fvzpk5XVBNFT/KW5BLN2kdNNOC96fc6BcB8VlrDKzlbIHJVVgSf2ewPcErshZXUQX6nfcX
1WASmwK4ixmJf8k736nSWBHwlLV4zKQwJ1PdPQ/GGInpyEjmaMaJ14lvz7g5+9RUlvIP/+tgiYbO
Ht06L9BQwbVnGXujNe9qVyn4yz48xgjkXHGcfpLxt/TO0iVSe6dPlw8KAaXlIDDiS0IyzIEQrGet
DQoQqeA22Oo7QgqENDYpDOkGM90XarpveWWW//g3k0x62jxYMZ/Yn++CLq7XOjtHyJ+wsj7FsoQ8
8ZUN/ABFKWy2eA31GlPFPsiPNKX9MJ5X5mhQzCmyTL1ewk/4cVXUY74MQ+59MT9+on4YeiJNJEPi
hWsyu03gOz7gb1Cw9mXz8m2H0bXhAY4JDYR84PdV77LS4eFZXJ6eQl+ODPmiPawHbdQuU8Zponz8
QtamYSmSNQVqDwH+5WMe6WL8qV23O6LTm4wT2/bb+ECy+Ujj86jF12iHl6Ka6AL8eLhEXrj5uAcK
p4bs47EPN7oBMKUJVy5/hxgUcgd8gbTbj1n8rD6fbhVbfnuMWXuOU3hGklViORIs4kkMHNrZSO9V
muhxLefVJnjLovM1LkpZV/7FLLFyz3cO32WwmC8ja5/ERQb3CwkQtXxUbTtoWT2CZOgW11JDnzLi
x7QYCLd6fL8Ek+8kHE2Ga379LsmNv8PD2aols71AD0zWD3zqWpAP+5AFJaKe1glukl1Fo9QQBLA0
IzWUuOcVByPkzNO2dcuxM69RlNJom3zM6lNrAqtyh6t4GKwKvyzlvvXRoPBI8P20/tW8cNzK9ZKT
kq6ewtQQwWDoz3CUxRnWlO1FvKFqkYKg3ruG03m5r4+B/HU3ZEgK+iAODQ8FPQx74fMD4DMnBu7N
2pzMTn7+l6y+RVy0t7z/lVN8YaFLk0FmtOLGy0E3QBE/1tXoao6+8u0+y9IhUiTuuOrRPZGjpcLe
V/mzqmrqASHps7JrHIRTMC8g7Id/mUwM3SIgL/DwwvNEDRc5K7EPuLCtXVfwYgwNN6s1BvDJR4og
cGBRyqzXlEUOZa5bYSlxpEX/6zBPN7DWpJStPyVFf3suup2mNEICHhyAXesvVpjzVIWzj2uhR5fb
x3IBp7HD6oH5gwaEPbKOJ0KaWhiPp8Zg+bDVESJerqLKOjEozSBKrf0WYWB33i8wnqyefTxBC1kZ
JY5DgRLfpoKusWZ8csPfZFfP1zIpTsH97O+PZmIEMbzDRHnOub5l5+XFFerDGU5XA3Xe2ToGZqRL
g4w54H+JClrm0hO2QYy2Lh49AyBrVk6oRBvE8/AtwosSiyWGW0CEMxiMTu3osyFSgPXulSMnWWDI
+PQeSbrAYwMH+37iwLpsfnrO5fItbhGm5wVSvXXymZxYodLw+kSmAKDvccg75DrknD0eioJD43xM
/2jeyJW2F53PrU88fcF4I5ExMjtyhRDfMeM9UX/pI91L4fGiKf+/DzKET1WnJ0X7LXoiKaxDJUVz
zdhAAWQzqy2XmKvJLlLYNIDyxGRlqNeUVF8Vbrl//yYP5CNOv8VoVW/VAb21BhTGKcq6nU7ldAmG
W9IPF28gcDm7RqBZdSvOs3wS3yDJA1WrqAbK3b79km+p2ybk8nc6Iiq2wMAaLJXPcrb54zAY75wd
mtAk24DFUEzNffalEo3ngTvlUxB7JkJnwq8zKvZGod1iGVQwun0tqFGXHsZl0Nk58Wpbaaqjbdl5
fMz36fEFnhTvY54LvZKeKbUJv5g6c1waYeBmlsO0HaoBm0SazyNPgejWzaRr7C9EiU/uvxOyGHD6
ACJ55LhQItraM9pJP8y4FrKWq6Zi3dgXcUKptaWtvfm5DDICY1NXNOyDeoLabKYEyqNhPiV6deXy
NACHb5dJvglrGM3pCmDHSgTFgclnL6ef3N9EXJ6Vx5VQt7/Mq2gnAdKnE+qfz/EL8oQrKI1QM08A
mbyH6kDRVSO12cVR4N1LsRfBCc44gSkRVsVJBUH43Esj3DSeAgiZ3cFML/Qln6ozB1hqlHZdV3On
zkRTGWOq1+gzAweVFXpZaljibMXqRzR214CEGte514MRaO1UYrP3MP6WfLqAfUkJY+aDzExUPB6b
JYq8bFbOFDM27AtOTtERYQXARz7asMFfl8e3jdFIOrGlkF6RjIva//kVQrdR2yTgtr5u+5ncMDda
hCt/iybZ5IeP958C6DYmyLcLSBNK6o5EOj25JmNLkn4EINo2HY2pb+s44bQ1C72EmluskKkgle4J
4BZCzZow8l3e7Q6xAh210JkHFtTR6Pyu6OLhY/3BEhakiaZaz3lYeuJfWYIrLrjUMrU91WjwjxPs
J+8iMPlx2zeV1hBNdy2GkhyDymJwhnl4bkgf4DacL7QWcEHhSjeiIqtLJjt2ymlihDk85jttsBX3
oJY0sZiDDD296qRrQiYd7vTba/SWxtAuN+cwaNPDVbun3+C2LP74iql2Zs7HDlUPwzlVMwyQQ8vH
0I/0kPwa5YeVNEP/Wk4Fon1hsfyeqp//OhH41rANFkaEqSBzgfyCO06o6Bs9G6lAa/Iec7xogfeQ
iQJe2tEpoSvdD2Xrg6Z4pUDnvtimAHwN8mBlSlfX9NPuZymfEW+mPfYo+GXr/atC2+f3Z6debVrn
+X+VGxFE55Esc3FM8575C613PpxicI+Nk/87rdnuLjTbF05SPGWDpYQ3UTtixo+XAxayoIsb2Yd7
7VYNOdCpu61lW209LoJNubZAMXRAtPmWb/YZ8lLUneU3SgERVDOJGkOIgTrfHOMgTU2l9KuOimdj
sWmEb/foyNlMOGIEKIavBLNVySO1Xiu4gJn4kJRacNQdiCe/FJbNs2gVrb+yBNw3EwR2sYODn1Sc
N4u5aj5qtd6aA8VY3UjuXfeUXkTm5+cXqUiUf2mDAFc2D1zs3s9wGScvOHKuhRgKhPNk8EXpikqc
7wUzOgXBIor9v7W8NBEO5YlUSny7w2wWnB78gehj+Z1vwC4pZkC3fJUTKTy0biIrInc2krmERZCo
TxtSzQCisw7EnJAVc0Eiy3WSmeFHGUOdWT2ibaP1PlJj/QP740neLyA334HBoD14XtwwEpXbXzQu
AGssl0x5sApP8nAz73CvPArziGqIQc2ZVZfx2FX9QA9gieyuAr3ZUazELR3WD8s3+16FGWs2++R/
HtYps+nZc/KK4MwwBNe4vVoQdjG42KkSi8j6yNaD3qqCh2jzNmRwH+wk99iqnFZcxxI6ETPIT3mJ
fn9wVeLpq2XXYsMzPYSxDZhhOorfA8/RTBeLYBaLTSp6QOh0rZ9Q+sScdzJFArJ4lJvmauS26n9H
da2Udlssbsi2fIM7hJUfyJt5etC5mJlhtvprVd+HiuMimhgO7V3hrivoTJ5kvmc1Z9IILRnOajX+
tPyj4/TgkF0lCXigTOWh1db0fsZ25YLnwtDiiWG3EDSLnXyR0pMQISS1jamkmhebXRYyLoqjwqWV
KhNLMyNOyEOhPeOhbIRTCoIqnBw9Nh58gZNY7qmGON4czCqnfRhM/dC0B2Whnh442U5/PmWw6Oxp
l5GeX5pHHhHETwsLCn3Gily1VDZefAq/oORnsVuW5uBV79dlHFWovYrUDA76FH34sqlX964UIMTz
L/NBY2qGI2aamTd+FwAycqc0YHKCzRDgJ+FbxJaL3ynUvtX+i+7JIWHQzkfMzZ/BlLLNjCFE0Kjl
xdmX8xOoB/DUzTKE5th++1D8x6li6+0DF9GuZt/1R34hTVDOzfmIAaZK6oqB6j8yVumq4+R1Mp6K
JbQk9KWQKS50NdAfoOOjIWYJSv1pOD02w0fhWvFX0hq8fNwtZH7SBhdO3Hh6oryMmh/V/NX0PEsb
g5uhSk5+yNNiEkATsjaiQkYvC1haMK3NI7Suc2+dtq5K2nar+HS3JH3TVEMlPm2WYLNypegpTzMt
vs44+2Brudh513TmRO70RZ9M6e46OfppkwFtVSmDsWcAfMG7wK3WhPIXRH5swnTk2CZvQeXEBM3x
NQx/GgjlLZXpyM2bYGbeaLR1y0EpqKHXQAUrYikLMBS3XFvvfpMZ3kHCxbzZMCvsvm/X46t6j2eu
RsDgQiaVbVy7TkvIH36VuaJJpukRN/HFt60/Sm6HszHGerxRySuRLngRcYve3OIrIy2prt/pzpg4
/oCOetdQ0UgCb7QZRwOU4mygDNohAvdZKrRr4W9pf8/H9BEtCBTyWCEdhxXHna4uH70h9KFxkD8v
GRVt+NbMdVdhX9xCBurOKmEV4UN2Fu+dr509iJYqZobEhlk4DxQNRmT7pGECaymdK0cyWMRuzub7
qHOjMKDK9PA4OC5U/V8qCPh+7o4mSntBExWRpDnDp/djkkVR+PRBt3///Dx0xJa5zVJynUXh1AMR
az7xDb9Rix1HO/4/MuXD27FbU2vynPBSam9qUE+BVkV4V1zKtw7K5m5ndcd9akfkoQB2X8BsXM0H
gvgnjggfenXqpXmkoFbFKJxCRh4TgFaYlN4OA4VVRHV9BWxYK+fjWYXq0hL3XUzn2dLlXiJao/dn
m5H6RY1eWHX2bZv55v4q/hwzBQRwVMLYJi0O6DKDUXRsgHusGPA0yySOCPhrtU6p/prQYb4VwYKk
hU7QR9AuU0lZ5WlSJKpo4/kLQOTX8Xy5YCBTtt/d0M/GVznOC0V7DkrMtIdPOpyceq7xfzAM1drB
/cqmWtHwC2Kqpk9G3+eFrt+C12k7eiZ8mWV+cdt83GYo8n+X7Y/EzlX9MpasPbhm608oN8nq9DMv
aSWczdK2f1Lf0PCLQ5GNdUJgn5heXq5+IaMmjEN9BG4bijed3dHJYUqNrSvmtzM9013QZ8miT2e5
PnufgnDygEAFjr3voeIvEzehRsH+MJFgeLPg8X8851FRvt9lAb6kjjnzuusOIPakqp3+/nREHm5y
M8h/neDAbPIhV71HopdVoniYVuTfRyPEzp4VEZYldQ6FeJkoc0SzmmkNLZd2BeD1lUFtGeiWpzGg
kDHkxvbeJbGzMOcKTFS0UvVLgzOh4BM8o6qWXW+f0MRXVXZR74rLNZPiT9QsxWiqgUYqsR3odvkL
XgDaDP2AQ/hyPLftJgb206S0Jxpk01isqZIHJ84r2XiVdeGdWBXQQh6zbiAj/0LOzm/Ss/SIP9Ml
tP7bDuu3uFuH6r0OY94+8sbPaRxg6RyOOYWQelXce2Csv5XWKVLV8WxxT4cxFEBzDMNxZIbb+K1i
Jh2hFo0qzQ8uyo7AIgqQBZgQVba0p3vrqZdeLgP/289HLunGqgWodtHzEcZRlseSOjGGY0VTd+OM
6guK+UMjzbLZAXd+kcH09PZHgGVplzZq/VglFu6j2Hczoh7ua5+pvAIywn+nYLi9Cbcxv8wTbpJN
Kly5RFcZzbzPzA/8woweSRa6Ty8e36ayu8FqnzUralfHdkI++UaEKGhUS1HwSyEzJTbYZ3njTuur
AaMeQr5ffEB3aRU+2Gb0PvLcyQFf8s3kz1KjNB5Dja3+fuduEyjMUsobM8z0f6fDJD++gP1IAcqT
LxyfUlgKfbp1S2bOg6/uBAUno+yNuyQXa8wnoQFo132vIi2QY6jbI5Fj6I7N6P3vnSFjRHz/Rfnm
q7JPLV8nJADM/iAy+K7ImabCZBwb3Yiqp76syUBIfOwDCV9paxxNz/qj6KlULC50VZTSQsDKvMiZ
wHrhKrnhqVznK5ryoBqV2daRG7M6t7VJlJqzslSYGi9UfxJftWF8Ie8CrFX1eCR+GdufQbT/0ADC
r1UG8fNuAZoveQHZnHcz/0cYS4IWFejX0JpVpov4QUntJ9MFj68jvCDZPE+RBbhmZgGEwHx1PqsR
MOR+HdTbTavuojCmE58qCEGExHW/jFy7CbdEmr1xuMqFzMEE7xduyv36gaxBn/KIpYJmN/f5lmyU
yrz2yPXSV9g4gOwz3OfIS8mOG5r8oNlIe/LypRGs4YMb/Fe+62QJseF3Z6/F2Aro+C4mTKReWnnT
jyV7/KLrQ101rXBbuSZZYu2BkVXIrBdlR5PASccMEXaqX2+OBE4cJyEA4GHlqPTAOzmdu1CZl4TZ
bE5UnTfSg4E32qcYZS1qg+JjhyowgfN921r+EaBbDGQ1wsutj1w6EES0YKmCLZbhkKBmakJUxjfo
/JiklYUdF/NaBBsz6BYI/XLxFR50UzJVt2AXHRvIquTtRv/TqpsGQPf2fnOTDQ7ZeUPif1H9s7pz
hMy9J1rzEgYe+DiEdnEpQZw33Ddm1zByGPfgodRNr5A0Iyea4Q7oZ6TdVFTWc8VRAChjVHA0nRZA
qYZmzL0AYbkD0zsyw+BJuKF6LXzApkjs0Bur1ftlRbY/Fkt+bxkSCSLTgM/tajt/jwJvrNirEger
w3WIrVDbRj4dbfbqSWaFym0IhvjvM+KkkMOVuwMyhR/ExOfS3ASaTNY1OtsljXmlzv7wW+arANB+
Mz2PTIzxRinp27ikyJLJb8Zwh66IqksR+r24YgWq/lfH0MQHcxafeOH50fGwLZ09Bq5etxWUlrRq
G00jn4D+4KLdUAj4fvNJSdRU5Iex5To1Ce3O0+wFGePMUCtFhN1Piqct2hz6uNYWLrCndkMXT70v
9tHaF4TXarvJ5oj53VZYS/hZIYk/ZzFi+XBfv+u035+CJZIBZg8oRTN/mNpheovZOpoDTL9Jv9Wd
V6wKob/OvgyfJ5/xKHiadbU0AWBkQSI/a5PKwQVykgsBjxTh2+MbuU/y7sbP896kh/A0ERHFtH2f
bl7ZyaF03KRTp8YZKBxDH1v3pALqmWhI5ktwOdiK4AKg5/fKBW3jCGsTN5uqKXZ85JHjWy821RzD
ky66Ax7lj15i9gDg9JHh2QwNb++z7Ll+UnmiTS5AGPkxVje4rjL/l9FcIsljCpEc1A/S0rpZR5yi
0y6S6imuJP4Ygtv47DFOYDYyGDnq98xPARBai2A2EEaSFq43/Vk+2hB0ze71Ru+6HGsnOM0c35L7
VkJgy5xKrk5fNseGm5/eF7YpF/2UWPumFZo/nMJl+yN+u5E6zahCiscGOZ1cLQZCnmr4jk6YwTV8
nELlgGXUV3aJc+HgA3S8STpSiTh/WUFVwdmE5gQyFeOAormmPjI8+aZia4EzR2gJU+Qg9uV1kPM8
YCK8fXmwcZtmNbrJ31+9OJVBI9mHIRdZkDG0xMVZdeEQB46Qt7ahm5B4xGeq9+YJbWduX/JAKCVW
e4XTxNfEsFhWX8SchY89F1ng3poSS7jVi69eGlxiRGJVXJRMgXIMmA1lGjns6Fe0lMi3Qu3KqMHc
M4UYfZSd6pFuMhhfzD00iTKLubTk5cDstfLQpgnoQeC0gD3zFUdjMWDTz7kOUbNBT14EJFUtfai9
kxZ82+OHzv0TQXnHMsHS7sbMZC6dI00yR9oMrdc+A2xv3x36VMTIo+qnVXkXXN+w1a45xFtySVna
aixlgXr7X8A3ti/eCZPA26FA7EERH/g0eCDPRtUT7sORW0nhC9fyxyP2XdviMAEQF3co1iwoixaG
4vBtn+Ih9bRHj34AGYBezNMYFqMh7x3wf0Ao2RpdOtRGZAyfSsvWK6mdcJnBJ9Ondpy8Y+/BB+1D
q2o52gkgcaW46/UmmgCe1EUoI5JQ5+0qbzZEGfgc719G+DuWwf84LCRWfG/JCAU/8Pc5BOvUYkfr
1iNCJBTFIuvwdBqrQPpksuOv57BRK+thSOBgHv3AhZrebTfDEvRV5rJTYALuLQsACo+xyIcVMXml
5qyOl0G377lILCRBu/UJ3FlOyODO3qbMyRH0GMiNo/AxpQiXaMwKX2e4yPomTr6yrGqni3RCx/Ns
HPWEx3UcBkDtyCWTbz9/oHmUS53f7t1pVL1iFBSrqfYjb5TCwm1uIByGwGPuX+3fo6LW9ZGW9FjL
2lRcDXYsXasWRZIMUviB0hNo6oMOOZMTayRyIcrJtgb4gdraO8qXsqhbzSZzthkiV1YaqQwZyOA+
qFN1MDEeT5MDHTpHMX90kSiY+LLi+a+NYPh4WIGWG1PiikypWkYab3wHKuAbQPdOvzY7Z54hPYpq
nq3AhOJF23A9rlE3uv3IC8xDVQCJ7K+1AbQXI8v2CxVaqs82l+Fnb2GqYz5KDNdMcWmn0DTxdIeh
NYRc7f+o+aBhm/QP/LZcJZb7K/XzYdWmlHgNrxGUi1oTeORKQ/iLrFnugdehi1y9+Pkj1RQuWvYf
AkUN92hCr2B00k0sgYC31pS1g5WkTuN03PUF66pq19lk5Yx97cqy81QMYDGPWN3Yv/SIo7vXt1W7
Cprp60Iv6mRdhkdduNrem2xKvOZNcgKJNF+w5Tle0qtptjMbQYq/mrUbpKt+KfX1p2haESz3TDcv
T0cY9ozGafNijNx22GiDB0wArs5HFPHF6bGXNCpSx3MF0WSDIpPbhPGV7dAazGf/u7kzT7v5iRiR
LNRlTgF7DC5QTew8XqKMu2+3VdA4psfdWtgm0LfxfkMFkpiBrFoqV82FzLF1GVsEKBVPhbEG5iO1
ECCjVXjDQKHI2xMsmoF3zCFhXQkOV9v2ndr0net6OG4YoLjtn+N5dclLvVUetKgdkCSq7rJf3676
3ahvOlfEuizie06U9Od6SCMmyoZH2cCpRI4WK70hS7VeP5+9SRHlBVuesdKXHc+8QKM9IrigbE46
H6vyc9aVfcICQx+35vDfYW05wxynZ+CodQ0pggPbAMoycBNCqTps/H+WGuXiQ0zKIJ+0ShuqGcvR
K2KgJ3NPE6jYqw7spUGt6ETxaXDgjAOUhu0oA/DEHicq7kB1bw2rX0YKgyh3CcYJU6NUNFXHCFme
tf/sI0r8NqCgluOc7TqLfXHOXbyXJ4vamBAtgTxNZqMLyshEwaPRhWMVK9+hqzK2Jmr32GcTDAdu
7SDZfTH8hfAuOgwVijH1QhXRYF0VtMASyyi8wsfKL2XjcEufQE2iz6JdcM95XQveTEILEYnd8ezb
7nFFq4z3eggsXJd7/9nTomf99y9YKNaJQeAn8Bh2YFyR+leIKu/2XVsd49/Lp5Igxc3q2E0eiYgC
YxKD5ekCYNwCIIS+8d29kavGJ0mYRhj05JmC5/tAViuBms8kykAtFX5Qp1fzvErDSgOFORrTGW1f
gJSnLd8tXl8p+9uJCD1swUGXZmuSl9WLmiYitv/lomiGorBcrzyJZQNwezCgGKAzvKFxkBEC0old
aCQnTgbuHsYNPUcvTEM3yCCW/IzcWU09L7SuqEamRYW2Ra93SEXLQ0g7i0n4iN+BD12eykhO7oFq
D2Y4NeU2FZ5WlyDz5Zvhy+hFPwshpWJF9xDlO4g1ygzBKGxS964v3mNna7yZbRpNpOPmWRoLeLFf
IdS+HclXLLxeg5zGxzRIfYGFreP8/EKWhTZycQX1j8v9QQ9PVGtlHe+2pFdiAGfY5fh6OIEH3VJR
w/AkfUICApz8OM77RG2Wxh2k2XQqBNtgg8IQ48o+A7/3avHzQpN+YyS5IOrFkKLo8uFrTUNjIPPY
hQXex2FOBwIK6Sh3KPivS5k3saex6yjy8Vz8AO0H/DFrthtQG1zfqb4V/AYXFDiI38JpeJft4Eld
QEUEgJMfL9eZ2ULasdhfKQvMX9ZlwQLluMALgmw7mScYrO+el5UDFJr7gfBhm0pCEtw0XQuTw/NH
wRY84E2o1Y8BeU1MYPQOo6mlia7O5KylimKD+vN1OgCYXWfecszVG7EOzGUOy9RwuVvX7QWiPjI+
L4oQqLsrNTCHuvNjrxwf8xhkH3N5Kw5gX6reMpUS4KXgLyqj/xr37sH8DTpbVZYBBX6xzMg48tOu
0WgeGI6PMXxDUH+bIf7UtWqMbKqH8yHoOaMbUPqCQAriB4PigImn1WP3kmkWuFszJBMOQ0iAMdq1
uovZQ+7FTkl3rqAlTfPXD17SHryjbDKLieAm3wR7SwMDy4VUiHqy9RqqkgeWVc4hhcyUz/qQkEne
Q2g5nhQWjqL96du4FK5eo4jK65wm3x82B/5igY32GDP2NTLiZyesqjyZzrQpJTAclO2/FHPBAOZp
jHnjEZcm1yFa8YtBYUjMJSdZijjZz4enAHcPcp5BlXqAAfjbb02rxTkaqycqBsdS20O0zY2yKGr7
mU6NNzQm22MCMfwODeM4nwT/SuVVGA5y+TeNme60kMGbk3D/A00QiFJIShxhTyjWS1BIXsr4LYVb
VdwGqh0k8i6GYQsX+y0rR5YUZnbg4mD19j1/WL2U1c+OMnmvHsRQ720YxUG1Y5OABwj+E/ZlJah/
g17bm/Vuf7T2AjtL/mOYHO12BHmd1xniW6lhdb6xgYyDb4Vhb0heFBPGUI5cSxTkOem0PCC5/OL1
/XUKeYPNbqRxTLpqbhp0gWbirdQLHuSuDTprMx0I8mB/0KzjC19VyxEpf87hIwN/Mf0d+7P07VXx
bCBEiaFe0dXf6+7M07oTuFE3TyRM/7wyHQF4tot0ZYjMWmuB1QBRogbHiW7XKctEBgYAV/Uo2nSf
MXHeV9ebIUQsdkhgg9ZVWkyTcuNZjPbRWtixKeZ0AcWbwpqJWrJVmttFRUrjcVn2EeUG/KDcF3U0
6IjkXgQLt4HRC2I50SkTWJtgtRMCHCoEVajK7Nq9jr3+5CAxVnxpGyCc7jaNiQvJraYyImvaJXCU
WxL/5dR86uaHttjh03qtWKYo6k4IrWAb/1YRhXVloKaQnT1YMEKZWZ3wiCbENQjI2UU+g+yH8Hen
57MEw71tttnWU8jvL3AZRR8p57XuH/0+ZZdNLQ5ftvJNho/sgIcvWkiboaIy5k00Aqa5ehLVTQqt
lZTwUdDlnJrcojPeYdTlwy295mmYdeYX0eG/joDVZ7hxcKL1bY3Bud87Om0CQH6cOfG7wufQjmhU
qOnylfyLhIlqqphghCKbb0H2hgEGJMyTA4m6FDgiDYjI3BWt7GFkg7ZjssbnYOehoFG9mlJ/vtdP
7fEZ0OXvbyMUcdt0ANZjiz2hbIOEU9Akk5vwpDpUYmGXGI323YxDt7ZvEN3KpLiHpjk06LkCXxyt
eFzdKL7nWD5Uu7Wp+G0RvQ9Ey3A+rgCYxCfSc1LpyHu1vGzOYswqJtywA+L2+4MD9v0qefeT6rXl
LwWQkz9+4fvBaCQmEjEOk0XNhGbAM5D6nbvKeAg6fE0gwiRV8bGHS1iPjx/QEKWk5UToNs3i0Fmb
5+aRrPulkgHmP/dPq+nCRTOJwKoFrpXjklHRmf4msbJqpesipU6HE5Y0ky50RTgFCzYiA3RIIBaC
aKQNXkrITcNk8j1TSJLg5o8UHeeSZFn9H/CtTYIU3drP2LScX0c1lR1HihRtIsKFbfiMupWjY5xk
1JedF2Eiycn0wlAdN/zKV2fyzefmR/yk8BNMLAzy633wDcxir4sKmofp3uNcZPKEDu1PMTOagg3F
bG4SPFQ0brCd1sx2mhy7JWu4K6Hxz1tgiQZo3whCj3qaNcJ9u7CPY++V53cJmh9UEAt7yL1FbsQf
ODWmx/Sx7RDZcttAMz8tyLB7S80H45KqIQ9za6FZ+0irv395a8O/NZgkUgHdqYaE8+jrqs7d9DeF
6KnUnn2KfCJet1BRDXQlVYkJjb3Y1kuDzG0WQa5O4p2gL7bmVkTBzMjkOoUIBKomk2r8MO1dHJ5G
sJoRzFq+qOgHOG/6ekW1IOpLlGat/d0J8AgcunT4ZdAsC+y9J50I0DZTYnnO2QBAbl0PqA7yzgfv
mi93xVJzaOe/N58sA47Cry+1n4Z1/GpAA7/+7LpwvSpTLj2X2UwhXnyy7Z8k+blzs++qnTa2c3KF
5LygiPAR66So0jsCDoClL7Aj0bu10fdgcRmGVMBskJnnLADKrG7cwDw5JxPHkQRZv8u8g8pDpeiI
xzV48uRBbhPUUlpc6bvfD2cspvJNJ7fsa3C08hX8SUdKubdWyF17FaAf1xQnOrZKhWaoiWIV1ioj
MAic6qLWvCJX57cWrkR4iUjePb4xfgWHV+WYJny/xSgMPc389Wf+HwJvxjUnypKXxXhSHNEJCkxz
h64jEGRBoFkM8QIdJrd29hMTW9kz4sJS17Kbb2Xzr72T6dKUPBiTf11x964Ujk5O/6wnZ0YjiIJU
Vd0+0H7XjAWlUsCCorihkupRmNJZA1tXX3+Qz6I9cyWZe60ITgtCi2qRtku4q/WNyJ5GHuyzqYOs
8SRi5OEi22p7b3+bHHyTM8lw7nL20dHMIyECGCok2tl4QpB/V36S7WUfezrkbPnRuFOQtmAEJY1Q
vP7nMcFAYB0e+EJNfpFyRJPKeDgQ7TxKeQ9JWMV/SWv8lKOcvODZj3s1aoN9GM5FsJvFBY2hYCiV
uibxnD3urwPqRBhgCy1Vqyp+/OPb7ClPAx/dfwXUCXVnk6fCOw3QYx+P3gFVCfcWVkZ85a5PRS2a
Q0TROzi+7aHZlWk3Hkm9aST048g8j2GuQqG3/lMIiD1REtpWOAxXk4BzB1c9R/oPVNS0EmsAJJoe
8Of2x+egPbXJQO0+KphQRQpx0ioXqaNHXLOyjvk5L2gq/c86U9e8NXO5fdTxOHnzEDnBRt5K/K21
R2XWl6ifZuKAdj7syrl/JRYt0V9am67vU7D1fpoNRHqwZnJkGCfftySbigBPpsKNFYAu7udKY4s8
EAiuZvXqFWHjyl3DBqKUyaoMY0VxXHA2fcCOjNmTDS13uslzCLzrj30ePds/476us4zyJP799Qvh
oT5SpXVpscfjI/tuY3U7WL+OCDP4NWpKOmo/LvWjjKUDJRdxUo7cOTHWLbKDUhGPB4OzbGsjj56N
QgQGIdvQgVOpK2Eq97jlMzvwqksSJmQ1ePmnWQHcnvVWAJHs7R0to74tZCkMNO8wvee/udl0MV4Q
vmdnpCSWhM31TZ7t2Mb2PDjXDbipNhF7BbK9tkrb6h75/yahTLziWOtYgmHNIA+uzT9xewTxPa8a
V0Zbh8mJfokhlsaEYWPJHuOFM85t/RsMohYB5B5Ig3Bvn+mWeYraMdblOsFuU/h8UPHeghoSzsU/
XD0695y8kN9ov8T4/l4IgOS1tC+z9mFJn61URaYNXm94cpJPx7tDgq6MazuVSgO9QLN7EFEKOhUD
fuN+zBax5iD+v2F+L9TBDjsL3WByxBd/fQu9FE1AFnWad5lvDueoS37k17+oDIbS7lrwppTbx0zC
9rgVU03ZIePQXrW6Fxddgl2PkRYa4EjVVJ3fnH15dNF6XZifYuJ+FdNMxh9RXA1ijt9V1H6/19pd
y8zn4dACilnQln1oDH9n46esY7iAtBCEID3PptPweOaJlQCRZ79UgJZksU6GBh3rn5bvNma2o+bx
AakiWVkHi+d0igR5NKuNQojA8k8rE3Kes2V5suhmHbpQNEUtFd8b9kQ6rnTFV9qN5JrpIWPba1ak
w9nRPy8Pm0SvV7NCdn1wNNYtD/qMwVccTpcqkETaDAjc0OGU/W5u+Zo/pJa6a7zaSqmnPeT/TUMw
Z0JLkTrORCHBULIk0NyAyUPra/1J+iY5Fqz3nNYX+Tuj82A4Xpb+B1QpNPBEtlNFJtcv53Bx9Ks6
bDo4DpxcMDBgu5ngc3H56M5k+IHNFBIkgKP6xpv7nMB0jmPjTHVOeNPwOn4u+sLPPZZ9S8HBpxGN
dHKqEQIOAfhItKMzkXDxe/Km7IpQgTTOaDTL086Ow1xW73Q4q/6/o9r9dUFjU+WlIifNBxlBrt7h
SUfgOP4ZMNhv5vsEeJSpPWd9+mDARg1hL0Y2eImfKS96b37jpSfIdZhGnjqtY9Jyk2h29MdiN2kX
q3asI/h55wwv2gA/Ebs4wZ0nQJ8BrO7md7d3zzOkBdwr/RSDXpc/ADEoWax+3NiTXHWHl01+d0CX
gaFsFA7h0pHhQkB+C3Av4T/qiT6hA7sLV7HF9py9Sthg1+fdxgARyGAUeQbPRrp4hBQZ2ooaar50
qKLdgL5IkWuQCTRi3X+zaldBV/4LvVLm4Q0k8JALo4NPPHC2eVw9dZKkN/Xe9ByfK+DCfFYKV5My
JSuiEcBlx1MyjRlpaPB6n6rjk/ziE8uGdQEdI7P28JX/bpx1ws80ax6YyCsLMeKcxTXfcV0IQsOT
sQ3JP7xg+Nhmp8VwfvULzrwlYqgC+y3gtS/roFNEwCQY3dPq2/khpClgUes+Hn+F30Y5AEmhCf7h
xk6ULdwcyhhEDxxPEU+uahYwoLqzfLoQetBamzAWCoioTMUZXLA2ZQAYTxOILlnJir7or2skBNOs
JzpNkHDAumR/7GrVu9SmgY1uOpOHKZlhkw1UF7KjVO1Za2Gtw3TWMk5YDw3Zc48bimjQavuuUVT1
4iPllrFlrScIhBzhcWTgRnzs67Dhil+a2l0gmjam2H3M4E2t0VyQumSRI6Tv0i/t2C+OtfuHMppJ
Of8mPesh3Sv7dfGrDtR54+lLQL8u+CxGPwspYOVJ6byyEqvBwEvosoBhYIjhvYzuyeqp/h4yTbur
XoJ2vBECQPTnL99H2oV0s6Wz4kAxCycAvIDG7+xmEjpivOtW/47N78vjjnDXONDR0Xscbbn/lqGe
1VRln1I1W0UtTPRDGj1UISEj4/tkbGkuceVY2/dHEUgKLyPzwDPu0+kFR7POs1OZuz84FksXuy9F
H4VL1QCn6930rtcGFzXBTKh2cLocv+KYzoa82r1aLyTAdBeG8cs3vMi7ICyrtwOzaaZoy+NkMifh
izXGnHlQCKP0yYSSekQN9nk33DzUJlrBQfyAQerOqJm7GLx3z+P/dBD6/21h/uBBQRpd1mObLRWx
9sMSxm0mdPWFXvWLVbq7JKIEdDL064oPbzsd8m6oPcko25VXVWY65nxN+QguKlGwospfcDj/vNrK
xEImQ3apagcYDPqoLz9zLlwzE1KiUTna64GQac2v3PR3EYDnNiONTPLVlCF3klaXX/bcxMENknvs
NTdUqawcwxyl3lT6yqy5XnJw35ExFjeh8Kd9Sv+cjh4Kqi4eTXLRA9UqwmPyj9FiRbjZtL0sUjx9
SY04esGuVX3B5dxbVHVLpSS/EaLamn1vkQLreAEihupyigmbruqA1RPepwtTv39m+PUuAzRz8d2x
OahBgw6EdjOKZKVWlVBAIq6Xirgd8QuNw2pjU9MAFyLakCtzBNRvTQrz6kvC/oWMwcTZW86pml4q
nQj/lFkK9UCZsaMVQ6yc9pFaHa300Gr6KIVjTo4uACFz85vlbG2huYy1uIuGZsNAZcRsMY8SRmyK
CbXtig0RDLRCiHXqYs60bLpMhyCQKMYfis75qPfMNClRqtasd3qhApG3ZkiDXE3TsRUnweG2Yyma
cJ22+wEgL1XJVEni/NzkbqC6r8NHlgV6sIu+Ci/LwUIpsxrBUaPVYN8aL+YvjbNJRmx8wgR+gtEW
/8kI05Y4PTZ7DQXvMbzhxC6c0QpJCTbXah+o4PL3HVrFjir+SCD+qZm3vl95+5jNhgzMSzJQmntX
4igR7NCF+zOgGKHlLnWiALVKr9LD7z/m77fQMxEFCVsgWvfRcRJb3e/723+1Ak5ycZ/GM5ebsU/V
AfJhLfhTVlbPe2Rulvqo9MDfZJDFRoJ2GZV1ldlGDUik1GYw7k2v3XGR6Of68Rn1Rd40EzOBhZje
xeOt8Dx1yNBx38a42DwaOWpaoqzw/K3C/JPtZ8oGGQs60UwTOFv7h0uvpGa+JFnsaXu5uUjSvwrN
4G4WYuTpjHBfUpoNgEfXzHk/iPMqk2AGLxy/4zLGU2ll8g6xvxxvdNDQE35Zae7Fyrhig457T/Ug
jBh2184Vy8K6ohKEUOjnyNAHYpIICWdpH8Sn/LmdjPT7OJ+RvePtozS6WvKonhz9Ge9+Uavg9aqV
6qrlbM1wgVZ5PL84fZ7BCvZAduWTMPOxB0jEUEhUJtPKTmJTryjzFueNs+SWUk4WQ9rgkONhkmWI
sYHJezD9RswpBg0VPyC9XuelzB2kfOkJgtcDKTApFcIX4ShAABpTS8YdoQm++G1aYtkwTRVOmU41
THpg1VrpqOr1ZMlWtBI6EUwfoapT8GqRGNGFY3vOPQRiX3FcPdZ/3mHJqeYk0WrwyA4lSeldIhkb
kJooPhrrLzBigF7mAQZT5enYOXLVCSWMZSFun+t++OEp2QXm85h5crBkf+Qpg4q0+lK8FLuasJvn
2udRmdAg5kMpGUqM4lC8lTgWB3mK6K1/eD2KQTMn+dGAXQlyNpdWPkB+tiQziXU6HoXyw25owXmw
aDguem5Ib4n5tRvlBtpNOD1tbJwQ2eYPkJEjtnsoIqFKM7WKIn7Gb2gecmBsIzOrRqPdphS4UkMl
sQY6MWzW2Agw8d3wjM/rLod5Zb4uqZxHOoYKwXhyYJBOjdUcYFwxiCvzjuX6RtEYHCsuKw7rd1dd
F0jqDvcK+l0AhGPj4fIS2ldNbv2oKxhWzJWoW6wZTVAUyz/Y4GDTEiWG0iFuZ2fZVON74myE3i9i
IzT3HOPgSxv289qwXSXnk6a8OIwhbq110mhmhCDfSNilnA7cgWZBLoNBqXUTiW08TCOfjSelSqcu
PJPMU4o3P7k6l/gCDENDxywfg6z2S3y8bMsQc4yjlm2CncsAmY97CyKKP1yogVZTjtlR0dEvxw3q
+A5H+8vM2e4kV0nFoxY1c5LHwS0E10lLO/QJY18KDS0yaH4pBUsb+WLuPfXh9ea7F81XRoHC67Bb
9RMx4Qp/belSsd2tCcZQZ90TFWeMw7JGG4FgtnU9YCj/Wl9tHySWojz3tbdOoh5nf/3nPlytmupn
kMILLfwn0B5x+ighFsOtyEUl69DQZEwZcwsGSGLr1ujxhb/RVypIHZhINy86q8r8upDWMcVhZ6hB
71Ao3AaIfEaVHcZz1QaCSIKbovnB2+R43rcQjIlH/bEUt/W4EptudxAukhzNHmPp/1INpFM9y65u
i/hZRrDvoG4ev/XeSMMkrMVDgTLTj4qw3ORcHnf6hdRlvVQF4tCKlI9kcJjjabq/wxjTue0wQgNf
2DVXzsDkzqg/8zlk8mAGK1/6t3EKYixGKh4uDE+dsQsOUeCPEafpmFo0GNeD0plCZ8IzABncYIVK
tRycS+zMeKcrJSSlaRrgLZcKsCnKMbpdfv4uZ1vJWn/RFOQLdTy6hQf5YfKRqiCt83kaMlDGg0iY
/AqsDuIR6byB6xqtsf/TRqYmYpnb+j5ZbhuVJLvF34kdaici1d/t0i91ORUDZ3JinjrK4hREsoZ/
KKXYhLel52eAkurPXeF8NNmgDk8dKovaAVWoXijxZz5+led9m09jQ0kUzxAP57E5zE+FvCuzrksh
ilradq1YqW2PA5dqBJiPiRmuDLMPaTtPJKB2uLfjXzC79EvpVJHkFAdw1yASi1MIEBHr9CC9zMZY
HL8FO+bz9SXcSj8x/XMewxkRoHbmBUuruxtwaKB37wzHlkdvsbSgFbQeJ5VFW/RpByIGOHq3X0aY
9W/5qhMlvlcou8LM+6Y2wgSazB/TtfzitR0JqKzB0z2KME7grDlYKkvk48r9gL2BfqUuziZoBWFt
Pdev6U7HDo+Bp2mMeAe6bRjMZNgFVzq6KLpLV1+mVuvqqLg2+aMBRfigALlWTg4n35wtekFkEeLR
jbPqLCw5Xi81WDs8X7OT1Pq7He52ekDvVq3PQ05mir61qze44ky26Yfoq3IZfR6+0AWG+RmVDiwF
sYcghwapjUIro07k85+/M5tU7CW6JhiHCNIiPE0U3eM735tHL7PM2w03hLyAtbxnLChrwG5gOLPB
gdtYNL/opG1sHoF/R/97XdAeMUZcR/oyfA9BjKechQc+RvLKmrhoE6YqLIa2DVSb1FOU5noTdgVu
Lhz8Fo4RajB47IsQ7uoiR0aiZgPBukVfFW+3PB1pZDlCpUZkf4Lr7E2WXGZfCOtpQnN3Kmlrhgi7
wwpp7gWJy4VwjhBhigEsMcST84/49HK4hV/a4zuFoKXLsVjmdmFTbI4qfTkRukcdcTytpxEhwdNV
ru0W/Y3OWcWMR3oX9nzM7N7cebvGvLBmfbRLw3rvdIo5U4WMcYQP7PJsh7yC4x49+PpDhJrXvCt+
mDJskGUYGtthcnipBKx4aShLXyl30gFhSeQCdJr+MNbehUGL0NMpAdkVRqCh+wb/9lp2h8hmSLLe
gUdj668hhwDWz/gEHfX2dwaSgEMvS0Oe2d067TGoCuFR9XDFPwDIuVX34+MKBJqiCBw6lMxy8ArY
qU//Z0QuzG64XPnihaRMQ+2iHKl0f1ysF1tiA2diHqIoirKteTFaZ9BFm2sl5j8HFdYplVnMlbTr
DSNMbNiO8qIPErQIV59vjNdiG/GhB8bljyK7d44m/Or/ykvJYHOn7Ly+tCJ4YKXmpZFzn0cyE3ao
j0ACXbkyU5dOzeL8Hj44QKVpVeABDC6uITxMBCFbKm8MvoVhZKZbcZeqah7Kc77Wf9JXSLR7pLe3
ZMdiKAg2hHHKJQ/4s+oD7iw9N+q3PUE+NVbZzNIcma1NObf80I3kXn08mu/Y/r4bERDjIBBXB+wt
Z5Ke287RdKnWhPwLEYBkXctRFpcWZrRtbzKf3pZPq+TnZAe3gDd0t5B7VQ4FoFcWMOidrTQ3VB5u
FLNbNBGKp5Jd0SNxajq2mQBR+sQOeHXj53iTuEUNyjyP1yyF+HACZL5x5AOjryC9jF/syftgjdh3
rCuMCC8D/pF3cebFdpDoTCVps0YuK8nUYmUb6obTmREQlq/ARqPByTSi/RhapJknMM2lxjkAGNW7
/+Vh9rXARcUemlfWuJyeHjxIJm8Ci6OqK06awhKlyvxvn++oSeD1AjoL1SnwMVOHYkKQ7VLgEq77
d6vOOLNk+Rw4cl+S4+NugHwTTTFhG/OPTjNmG5MjtP8+ORqZWAFK53141WLFq6U6qeKyBOoa9DVA
0hZ6XbNadVI23+iEm5DsVRdAF5v1q+IrH+1XveUNxcMdoF6xkFFpAwJjyycWMmhcPl4DJipWA25l
5+dIvgCn2ZvXwJChpEH7nofIec7IpcJHvcRIVCVQcr5sk5w4F+AyQ5kj/FIdzSUuU1kuB+xmbQoS
FU87G3JrAwdo+udWLMKzciZTAC5BKNznrBMtzN5jZLAuWbV1is4i3jMYct72q0MAuHZF/jbAycOR
tcdGgIHwrFa5ZSaWTA1OVstCXr/RvzHFaYC0uY5kr7ltKBqnEFu7XTjrEYu7YT/fFb340+eCtVoK
1GWqcaQ5GGJisM+hCMfuMOGTP82HZCuWHmRSgwxHCqf1buH9glTi8mpsgWG2AVMheZ0wbwAOkqAN
SxNn15SpqC/WuqhRc59P54vZl9wlbiaRi8ldMCgnFP+fkenXKzuRpGCJE5nR+OYz1NLqEv+oNtJC
7Pom3rDnGpXQBYkHe44+5cGbyPJ+Pj5cxFDW8sSMV9BGr7XnRjXco7OwaYOgFEzRijzew6mCMpen
9LfL6E73s5cgDk7XPdFAgAySfNDFmq/JHM3FTziyAEDugAgXK0PoB6s89151P2zl5+7shCgk11pG
LP4C3xapyl/SY3yhvTndTvb/Enri5AraMacVpGiqn4qTRCT/ZKQu7ueHG40VmVufrKrrHtqHChVv
YrvxavXt/T3m/MMbMZlIeAbwVJUrmHAYkUnQX3MLocEOoZPR87sBVziU0+vh0MyhAEJvoqVfigRW
6IxT0ElVajUY0FgxASmVPzRLWzF0ZI7AT9CkofA4GP6FmQrV38cPGwe7ffRNSi/NUif5N563Zb8+
fk6JtyGLC1QE00SF9WSBEIxh5bb5/TWftJjejQ4TAq+qqyp1EEMQzrCr8SnEhXDmNRIarJNa3BE2
MRW7yuSAeGcB24F+2SAPnbZmUsJBXqFjzxLVQeWl0gPi4pSZKRqgEEspX1gREQO//W38tSWLco7W
g6E3TK+HD1RLbB37Z0Mkuo6h9hJCuqydEiu/xWlNH/dknIuatn8TghILxQu2ys0tBj9aSNsl0edJ
DHxmB3C85AwF5TPK3foYqA0vIeYEMmowGsYCs7NAY81QkgDui90QAAKvkoLrTdM0T3mJ/o/2CXTz
cT/yoItyyhhwRwrGKu6Ao7VEhcuqyYqxm6n55kxBDvWlHExy76UvtK2nZrwJ9r56PGdLiZP3tJ3p
C0cSNdzYRYbXrTWw7Jc42GpeONJFgtpzJqI1Snpx8GSLYPR5cLvz574kk2AGUQfURY1oZqqb4oFR
c2rk2QPLDlN6AjOh2Kr8hpn2G2sbVmTeamytZxJybdbMffkisKGPHEukJ/XZldFVE4baAg+vrdt1
uNAIeLG4PQhhFGlStl2veXbTHJnNXjC6OI0BopjVZGpkQ0OSgcYa48bcUsZ73R5Pqi0bV23pXLSR
AI3R3MtC0aqb7wgL4N1EKjQcQEsBws8BLeWO1+4VYmS4l4jXpXLsFFfo5qpHE0FaTNhgqIo+w90Z
mrdmlNLEa7OLKP87VumNETadFUGOY2r3Wl1YEXCDKoT1bWBAHM4EYhj5j0whTW0X19isvOl7WPGz
DQpT7JWEVHOsu/rpLfN4ADWnRMfKnmuJ7989aeLfQG1EJ6QIGRHu3Nvyk6npQF8p3+qWScQZijw5
+7x6VlNxEj+H6S1g6jMPu6Zctond2gl4tNcLjro9Odaykpi4wzvJofjhisO/JIcnbleci7Ytolzj
05SqTaPppECX7i1QRkCY0NQCXw11es0RJvG3UGF93pdOHTD8h4FeuO0NuLzX4YQ2x3cuZ3jolxCC
RilX4I+aWY/UnsaQfPRvWWXACReisYMSjMM7Mh7GICF/Y8cqrDyEMY0S3Zycy3A2QrJUiKP+bkWs
kZeZt7CKWR0WosNifW/A3C42I1SnsKHDEpz2r+VqksEkfdowfw3TlONLAqB0EUphpFLP5kCOEPsu
jgPDeB6da1FKjaKYg+PKcmMqwYL3EoU7MOJRetJsE/uI+cHEB9mb26WUltYrpOFKBCAEcHQMMF20
mAle6TFvE/u8dyTKpykUnajhAiNFDR07wlhJjFtl6jACVm7iZQqSyk0V1HvElsP/bQ9MUyGlriKm
ZZKpKOlhB8fWKGtw9Z5vfXjR7sugQhEuM2yYVcz8rEMuP4opeQW3a8MpZar6RYqKcKUX5RWFxFTq
eHCJk7IbwimKPfucKyvCVn9wi/suZiU0e2nOWWgC76Zx4XJzuTYb9dLBhteDa/BAIfMVrrU+dcwu
PItCjlCtZZQEGfzgFCtVfvYi9kXUhrierwMyn4RM+BYyxYba0Be79c4H2BorLg+SzRTEqIORq8mo
c1OElthPqcpLX8hTwPuIyqawxEiRWRHGtm4/3Nidx+9Eoaec0DbnuObBCMe70W+qs9CUE39z/0Ed
jUHpMsoqnktZxr4ueDXdDEkzZBN5LItvitjfsUOs6sMw7iErjmoW/3r6pwq9pwerdBFvsUVOv+q7
HXAWLV7JIdzig8yGp0cFa7dHGi4gBxb39osDfMTeemiWgJpJEnCCTaEVt/Mr7ppJ7dmHffVOeaKS
EtDvWp0xARLPPS3zBmlUun1Br4JIkkLLqh70VdJZhLFJHsm1/bDfy/5MR/4m4n2SiDAidTatilF3
q5jCdSin1Xmvk6sjzzmHeDlQibbjwJ52MrlZL2sx9k/xfUgI6n+3MQFNGzEmeQl6r/JHTx2K8/PM
io/WTLdjuE02xUboSUHKDEbLMhmBJhntAQsDhCql4OIf/4tIGNrRI7NxrU86MFEdRiF0tmBJzB0D
IMvQp//ja1hgHG5FEPm7aMklg8dZpvqxA3yuTveGie0wVE3kHvRqbYwS4fX9nmO8pUtHFc2OyJMx
deUyNjAmntC+VDw1L/UnbBhz+GUdRwMDcpIzOE/qNffvKM+5nwZYWNbMnk1kvZ0hgjhlzW+9Ntz5
DDkp7W6IAg+3E5pQF68IyfLOvrME8nlzK0EgMKJ3XNRw5oJJJh56lQ4+usdVJ5ZP/VHMmc49pdj0
W181hHm9YBHhDDgl/LDNQ8kU9lzM4XYbhTrKEJ7WvuLPYq2dqVqDB3quOiF9BMHWofTv1jGdAmFR
tg1nSnHPZGaWhuZHzJLhFBpTjUpKjPtDV3hbgmtvQ+Fl8SspBnuYZAlbtpc6OLeOWWumP7Puyxjr
d/GDxoq5s57kYP0FnMNAABmjI8LEGbdXj6a0sBrLLgTq8UaHoIid4LzYcuD+0fSlbGbL+gxqFeh5
E5G8EWUYT6G112cfGsemuqt3IVJQ/l3hkC4bVpxNq6RiRUFozYJAaOEj22ITMWZxnU7m4hZomQcd
/PD76LFoAIZlBobwBD9fbSGMdO4OH0m8ewJm3zpTmGeWSxzjzEsGjCHEc013Lmo7f3QABvIaqrCU
Fbd9gndaLDvoMzlewtlDljZJH/HrrpzWht2TbT/JMVo5Srx2EnQTqpaKiVGMgAKJ5Nqbhn/iyd5M
YElc1vrnHNBJSywZzKtYTgAVHWPMjhHVZJzlI9hKYMOG5g1TmARlRB5BNYxlSwgzSeGcyQ2/l8ha
87fb+Moq/O+1QH4Xpi9qeDUmqj0MpjDLT2rwmh3o1feIZYV5V2gH/NfCoFMpvPWii2TI4dJnFPpX
qDWmKZhnzT+6qcOOeeNbWcixm+tSuzzOdiNY7Rq9FtXuk+z9xkB4ktl1JbeEzPftCgtmF4CzrR5V
vlBnYAfneXHRnZhD+uR7lrMh5/yH6pX7NzTgih/p6LzopI4cP6irs8VX5nBoq9yUkEfcXbb93aXV
zh2hFOfK+bLk/o96FH/e8RuZSupbqldJ+FNVf77cW3V4sP7iixtBKAQXvA8QHK5Z9sBsmdfyPY7I
vyMictvZoZ/biMCAAucsdJNHKl+j1H+Bc/+76cyP5h+QNcln8Ie5cnHMKFMLOLpXkX0Y6F4fnWLT
dZM2JL5QDmXM9ztuxvoxH+P3K5007lG8aeytctLGvQo9iBcrbowfrD/2Ue3s5kkd3p6uxUN/dNlc
23N9qZUH2mAMJzEWiEn3bJSRNSBd5lmpGtZxpC3GySBU5qOhINfjvE0dmyYv3lhABZLiiVuuK7PA
W80/5nePvCXjqotAqcw7ejpzR3Ur47NHRpNPIKgspLW+qd94myX3u3ii2R+GIpDrZTGIgs9JcdtL
gYYuGZWRb6skamEpGwSsIWETgHj/Vpf/g2XJ/dcQcB0lqD1fDke4BSbip0PVVH/dNWZSamIxiNtc
zRX4G2haEZvHrNZVswCJprBy2RD+rIsDab5zgTA7pGoSYDlgeQusRKiDIgDyu0uEgTj3WRjOAHSJ
kND177EIYzE2QkLedlEPtPgzJdYALF/PWEdsp6DlDAvYbGgJK1WReMU6xrxUK73QQqtvrfffOz75
082cRN72ZnKH4pnX0JYfL4kFQkjOSdP2f/qM/KKybMQIyB5eDBwcuHAZrvtuR0u/tiJyDy1wJXTg
QMP/5VDWLATkrE1q9Ofy+8WeIu6ktX5wC9+hX+CEzPF42hZL2NkBCpMVFPrhXgtIOxl/dhCbIo4D
eHBoEZHP/ZWDtLkUjG1ofD3kaBEQMsxuK/xEN52BF+pd5WRdc4yQj9PEWHfqBXq6EH1+GASjNNO4
sBv6Ck+CwGSwVwGpJGeDQSblZ5CH6kr5EW/j2leldZJIpt7/gaQ3XaXzV50e3BsS7+dhLjdfzff7
JXcF2N1JthEZSuywIRRvOib/R4TIhqqT98tRKfr5M4XYhsbihN2pMbyc75z0zl7AzwqUj9lSTVCP
LRjk6HVKM5NGp4Y1o5gH3ZLeaAR9gavgFyxYbfJf5uNBJDaUVvijtgCLFJnmmbjH6u7McSseBxbs
oZ4vtwlM72VIktbIueVDKG6qoyPnnLJ+MdBQQWhiFwUKZovT65FvIAJwFJrHoMKpUba3yjXflSBw
BkQm5qugEqgKo+m1fUF+/cDMqmwp0RGR7djh1O3YsjHbA1QH37pO2M5ZDBzKX6myxjmGZ9BYVelo
AA6vKEaCpZbIaBa7knVYHEsq48Ve5sg4lsRXQWCPbUa+0W2u05vZ8pxYuQnADgcJs0Fah1TPf1t7
U6mCNKrQ0om/bmgiAeTyz/GYBeh5xySF3fM18GJC5Tbww/vQp/Qs5LakCE1LFqlwjTU6ZWdA/PNr
8SK+4H9Q23feBBrCZf43s22IV0Y/RLmT7MKkcLevpuxe7XbKEkBvh+HGmMEii0CPRoZo08CHWcYY
y01rNKWABDLQqUvxrrEM+2NG9adKu64Lp5UosuP5jGw76vRgVL6YiItQO/lUFu4FvuW5CEpk/N4N
Thzv1BpYxEAQHjavv8Za73jzQQUGIrf5sed88O9/gsi5O83xTsVSG6gI074AVL6pR2jM1ZwnF92v
BGll+lCRn2JGoS5QSx0OXbpqaqgWkH7klftccQ7u08gAJNOncdH2sEG90dKlDcWKhCrEv5o17a/T
yAbDP4iDWLC4JeJDeaF6lSgmqHrguD73/u26a0EPJ0LvKkRX9Evpe/0LqI6gKwKb+L89cikDnRow
XnYZTp+SEfbgL7exO+vNLJeCaMm6r6aFlfPbzkzWFtzBdm5loh2lqYDEEYFPsI9zx4LTXZgl4f6I
j7mveDHSBn8f8Fg3P2jsg+JjS6hSqkKw9dgNjX7RaM1CBl2TkLqLODkddKp8YgwVa78etemzE4T1
ZFzZ3uMEjbJs7ITP/vFvG+W6uRnc5GG15IVBEYaDMX6jOy+JacwpJTIuUfK0Ga3nRQelvqba5Gc/
IdO0jUaL2n6YDo+9APrwxTDVL6xnQmEspNfhPeQpuxtpLyB4JP8/NeXHEMznVt3dSB1weIyqiao8
HxdcQ/kgMViaHQawxMk7coaJ9Tt8puunhDYVr60M+pqX20D73MAlo07zdv7ssY0IZ7UZm1scRB/z
skgnUWucK3Hwn1uYnamVD2FpxF/EuWfkmjjBrXyKFam9n1dwMQNgB7zdRS4ug4foQBIoZojXIUJx
s1DokltGkmwltcOtRpweYUm/AQOM26Onb5/uJaMJMp3+a5b97rmtlqwVWZvHsFdY7VTmC9O5+ZeN
ogbWQsBqItA/iY4f5p9wmD2GzrXzEUIHM83npByOYrIeZQUUpFj4mAN1hbQvQ6G541byj/vmYZtv
sPT0FI51zxP9SUoNqlSG4kVYMFGdoIZ7ZnAUe4JsZsk557ysyYOg/a0iJSUZfYMDeq74fqT6IqCk
r1IyfrzWVFrfmAfMt5C1fjHz6KXdoO1x9oHOrPhm+2ImFcEeJP3Wjc2aFVRvtXFn79iI6MqbWmqX
6kIUJPekKDn468SlA6e0X54X2bwh6EFhUkAn0LOWc0fxqDXJai+AwbxKQ3ZpMXqpj0IK07Ys/uAG
a4pv+qfc0ZsY+KEeHIa/EwQbfDYIuVzs7ql8z+9s/ZB9E0xujEyR7O5rNoIesdxKfNPMKCETD74+
vaUctn3bN1imp5m5Gfrs2KoTb7/Uh5eP2I2i/De8vd2HZ2BJYWyp7rNBurg9SzsHUoKLK1m3wS6W
M7CV4JUJX1qwfTEYLaBcI1MFud0sOgca0j7dSxoMswYVCmjxImnoOk0hMOdthgssJvPsLu+HGJ67
DiLOVQUXPgxvlD8KHgT9PFtuQh1y711M/cuXgbjq9hXNQa8nkQ2YgIPH/9Jpe4tiTURYg5atcRv5
h5nACHyQEwVRi1peFEGGLZoXPqOYfgREx1jTC0tSWzT3i+pb3u84eJQAV2ahTKJvVE7YKNuYLUsC
nTxFsSgjdtWL+xim988hQbKaic8WYFtqZUdnu1l15NSpr/Mgm73bJZNODnkcKYTMmj0nz4ZYNKBD
Mn7EZXaAbQwgjnqoNK/OF7OMszaH3Xz9JlgFN1bqHKEBT4/mtqedKkkgaGsLuB912CySD2JDF6Mb
Aac6/n08ELOEVkueZ8U05OcJEtpbgNEGlsEU2xsrm2kPm9kyKKpzv/VXzc6RdfkZcwK0rC1KmSFt
OvLz/y9vctBSOLx3vZiBBZGgVZ1C01yfYRhzgZbmkVYYLfM5oF0LrJUaLdq5FNFkKNM/GUNeipdv
3WfEgYnLoksaQF+lzKNdP52ott1vLheCOEzwu0RtZHffNG/3MKEwIsZ+WUIqdp4zGxFGYaPykkoL
d8HyTHVo5tOTAQ8obCe26faL6tOdWH3QfEUzoSRx71hxlNaKuhmgPWCgo4TzdCL92Jvjl7nBBaav
hwt5cQwSO2TZrSL4nF3/+PZ0WQCDMYIxf9qKB1nk4FZzWbWWsV5GZtsLqb318j+quWetwTa4jB2t
jEGUSaQZjl6n6x0iJC5LkUVdJ8I+MkLTshYW9V2VC+vJP8w7g4jp5L6tclpo2FTttpLvDrRZAHUN
dBiMMDZB1yZh3u265wCBdodX92kXj1DqP9fxmgZTFF5FrGoo02j3PbqcS9kHgyO+Vzt7jjJzfPrM
X/buyxl7VsPMjLdszatsYBkItcGxin/b1Uzw31EsJtxMhQ339lqilBYKKLRD5oVL+uQvQ3vmYEul
pm7krxL/Uqu3YQ8EYn82QkB71/XRtZH3k1/hoZqg4Ynm0ni/VRoEzNpzh1gAfGEIlzHiOexASspB
JvdhB+wJ4e11zGazRAC7Ob126I3J2OWJa6g2+AjvLAHTDzsxwG90Ap8Hl4YVyJuAZ6nBrOIcREVM
hfJAWH7HNiJVa8LuUTKcL/oId7BshVLK3NpzSOZAnupBxzRcDGlSG30cveCCI8EVyVDnHWTtFcuv
5NfXc+DE3wIbcQ+HzmVcNXIus1o1FE1XsHZCcOSbl5ECfTS9zUZthLJv0SM078cYtST1x7PYqo7X
zenBl79ZVoU04Adtd3XULjEufOgQlnB4B50nXo/kEJrFlDw6fQ82wUxb5zFFYmpKdIisitri7vOd
BFHcYflLYknoJn7cKlK8GMn0osorATEtur/54ZeWg4hcygAVAWQflJMPosbrvwEjEgdadWD6evmt
+ZC+Cjq0SEYCkbptMCpzzVpJn5EMfs9pXIiA1Zz8q5nnp2WatSXY1v+TrPaCH1P36K/+Ij4O1rtD
aHhWAl46VALmB471M2SydH2oVYPgXMtj/OG/M6s1HzFJd95vKHGKU8Ie5bP6kPS3WE6I0mATYhCr
roOrP1OjMrAlGWo+FkN8qlRvnYHXSivXYqbTA5WmY+yssfYwLQn6YDM3vy10fAFWQn7zxnscwrbR
tisYuf6Zc8PW+OVqQUGFkohrZkk/LcrZdY3w7dwc3hn9pCcOb8MV93aVpMM+Nez76q5dQJD9fg+J
IKwu0VeNCi9nG1m1km1ynHXdnPGIn68uT8Ke6mgOqphb/t7G+99/MzEgIg2DPIoUqsjPYTZP5j4N
paDiYPabsDtyE2aJrXFiW7DA9QrNdJ8mGk98v1ZxNgA0u6gid7SLrAoRSQ3/jtx/POdk7F3JqoCT
E/SX4UoYqQ3QpaMC/Myq0TqwpTG9xHrIT/ZUmgxf35c802MkrSKM+bqmFzZpVnoF+xyJi9owILcE
SI6PZ6SuznDoDtK+SIWhHnZstumIQtbkrAc6GGLRHNfzEZoE10cDX14oaVYIMo+QRIzcxmU0CgVp
wl41NS4VCd+o1GZmwDEGX0dkECAQ8lX5sQ+gXaKouTd3CS59y35c/TQ0HF5NpBZBHt/vCJ8kBNg1
SaBAXlw7qU9JmwfmZgpj6vt/tZRYnGVkUBo8pfS9p3wp4A3uroY2iWZjHRJiQr7pdSmVDxo3eyif
DxB9a07UGn3FQ2ieSHLrursBrM4cNYdvg65wGP9W4CZNeomwiqXlD2jkaxSeURd/G4+IHUTBllCU
lfA9nkr3T+RYzhYySLy0tRsHnSMr2Cbbs9IEzDTWHJnyH2tW/ul/FZcdqLPNo73PDvXFQaAVhRsW
yrsMlsHNqEyE8QfvKUtYU2ugR7VZ9OX/IIDIqjMtUe4KtKPlKNZJ69DlSClAF6vCd5QcGsz0kSGy
HHIh0pdDBIHEmPWe1vGBimdFX44jc6CVBKqBzOhVtA+J5P8hWeM3UylY0dvIrYri9wtCMjwQc/c0
A4/dKFhc3hVklRBxwkjF7LPFJoWnosyzQXmnrYKIkfc5W3gdJRr7Js3DLRlOQ40z72AeDC3PYv+S
BBJk0WEJE1ylkmFHZPQuM82+k8Dy7D+p6J1mpHB+HBBLYdlfudC5NjMhVbe3yoB8bANfKe7SLVcL
OdiIiboECUFxR3+KQofkf3XSSCWVZba/1gPoEai+kZ6YuulTnVAk4oq8mLl8TAoAENdmHE/MqxBa
ukd1NQrc4jkBKyojfsqW8KyRqSIW+EgV9C6RZILNWNxf4IKOonuEs0Veeahmk92qZ9XZR1ym6M9M
zvBfhc0KIGTcjRDTqZI1oAjZyHcQ1QGHGmIYD5C/827bpjd7zubr06fP0E5ai8AY+WwxGGeCRf83
t/5ofoYFV2kmzuDxx7NyH4Ev9zlDSM7/LbTjn3paku/16iOL8ZtHflV4RwVlAn91n+no1/zEO9va
azeUVtwCtz6r2Sba6G+5JYPoABV4FpK/2OxTraJFVGjvtyJbVBpKILQJkZI9gcKkCWfZ5GiulwBJ
1O8ZwWSj9SVUgbjWQlWbdKHfVzG2n+lrp41tMiAp+I2C+IjlvxBa1n5+pDe7YfR7Cif9oTJTE4EX
MXH/q7WlbDfMWmi0r++2Jkw7xy/CfjjevmGczV2v1Ryh7oKzqEsaOTPhCQgimud2VJWLNIyXFpDM
+RDcsFp195vs0VfGBZDKuyML8p1aB8WA2mThXj/lH9+2j73h73GrCKsM3ohc0bXyi+iONVe7mTCA
jMVzAbtXAYge/KPpIOEMY3kFk7eurYY1/R9CLUMIWC8XtZ6Bq4OXJMTgidrnSvXGWlqXrhf90O6K
ehSAt/6UZ4fcuE9gB2kS4ECNd88NmtLMlGHiv5jGDjP5YARq00yiXIYDrkNQqR2z59p2aRDuIkqF
tEtmt3qxaUia/eeXz9fnLhgJZGYoF0RHvZ6Wkz2auhLkBIGEuUhovbzhi9HWwLdms0d/JpOA3N2T
87ai1rFqZ1sgD7wIpHG1cip26+zZcuo8huLBKzx6q+QD6xLrxj3iCBQPkcFOZ9V1qj0JI2QFr4xt
0g9rd6NieA2wMlLqbyrelXG/+14FbJYlM/m7pEZ7MmekIxbpREIMcQ3E3YKXwTACwcDOArb/ibhO
H37SOnk83jCjnuiKyIG1go0alfqluVXmsDcpnh0VqDprN9Mv5yjYMyKJ9kamIUiWfhCut0c/en8e
JT5ZN0iZt7Jq88xkmAmcQYn1YU/kCKr8djTDw2NzqETYoV7PdUOeSHd0QEAMGVpOMeukBqTVzA9/
heMTDnKOB0M0fD9tmYkYnOtVdTCKM39HW+XGEIpEA+iwJpC8Q9gzJSF9FJ0dv7T3enm6np2rXrf7
ssPsqxTm3cuUBMpD3PDK9BKTN9sFu+UW8V/aQDBvDq3kjLkM6c88qCZXQSaOm+4cPJXmygzUSsC1
+lfMTxhNKpcQf0ytYoGTd8zKHckIJ7ori5kuPGL71QSieWp702Vzrf+J0J/aMc9e+cCw5/2qedUQ
wLCUS5pe/WnY5AOH7zvFQCby4VeC7m1Wr+BgcvG2jJkVJtsYF9baZgmzeBAL+xiGlB6FZRp6L5cn
/hsyhF3nBwVTBlj09JkXdW0e88ab/mpy0jrIA+CgKpdmWWy2HbCsn5cmwimIB0z4RCReH4WPIFVy
GRbAjERRLPyToWDBQCU85U/tmC3qs3hH2ffc5SYH6FbVVFUHXNySyrAFBrAw2jFoJK32s5D4NvY6
J8Eg5Khav0Lfl8B6edntEhw/LYTL0XCd8/+2j5mLlno8sOBx9azUw0HfxXG3EQB1j82bTJwtj6Tl
B4KEVFZUaI/ylPmKYKMFPliDNzD3FWhepcsa5aPBfLUjqrTQLk+hZtwmS5iBPgXY71RsQxWKW2fC
6+kimrq+rdR8D5XahkW8LvG6TDn9n+kadlgQmKAS+n0aEMBQKgwLjsI91sckpRyx2Gd9LtIRuAIj
iD8qsb4DRue07lXgJTEm6V4IXsI85WDAc16pjd9T9WOhpWQFlcfUZmidu1Q8wLDhLS1zXCZdTUEG
65bNoCptt55xeybkZRWJe+u43upRoSpBwKECUyZSg6fJUogQkFVJw4ZrRz+v/FF9ZVmTHSaonTjE
E0S1vKQJyxW70qehrcMVb4aYb2yFBTj6fSobq8EaklHJEHkMmxjUrDjX5AD9EfWjr4DRnJl2+yq4
SS7wqWP6L4PeIoufxaiZ448tmrBiJjFkOqMJ7oBgFqlgTicLMu/zPsRsoAGmi7PDfpjT4geAc6iJ
F0Ft3WHpp2YoxjLRVxNbdPnxmoJwMK2DH46TmiCL23XOPHSBugdh6jGFgnDINTaHTRwTUgojWI/y
g7etd3WFmyWP/O1uz3yMUf6pNYY/q1k1eVYtTgymlNJs5Yfwq5gjpVaWPs3kcdIeILN4NyYWhjje
8ZPcvoF2WF0d/IQcsifB0NMoBBp95XzXRWPt8wBTkXk+tajtfMqvkpnqxUICKXYONFPQtqAq5knW
Nzt5gXmZVOgeoDvGuE0AJHSDVeN2Z5ZHey0SFDkLjIePcJh0HFZypgDEK8fnODFP3YTmMrGaQfIc
HtU+wewrNSiCiWVhvHKGGMFKjFLxMZyzxzhqCVKg7ACcMLM+JcaUS8TIDEtI1yvS9eiTsP9LGi7r
9JRHxn8qhiQVgedM49y0J1CrrZbn6Q9xohF2B9ehw3zjUFifIZPJyH6KeraA8sw1fk1ASSpwJ9er
NWbN3zPU1U+g6GIZ+8HAgZu7eOaJaOxb9vu1oRaQuElMnn9MFwtCqFGhr1m5vir5fcNMTD+tgRp8
3mvq+fVTbAikEQZ7UhwZNBFwn4n91NnRvR1NnuP7tpZQ99SB20i7M+xulaU9FTbiouqBo6IyeZVk
zueLRv1Boq6qAUhaGgwCKY7Q0r3xpDQcn+bJXMnPPc5cGH5ryOWaSDKxJzcauIGo+dZB7I0dTGTJ
DzGKzBDSD9UiIjsgq9c57LsH1rg6UoGvQgMssHxtcss/hIgtJJO9CWJP7MGIxdhX3X9NiekSaBHk
Ir3fIEJQzh9LM1S0aLOsx5+UpNVEbcVm1MLrO20MiNM8mVH+n0fXnq9IUTXhn7cvSfvkEc3KZWwW
PZ69zEHplx8sK1yFpi3UJbBGQ66btV61x2d0vi6PxHPMMocV4eap1y8xgY6MjxXVb6WZQfcR/OlT
HsnGucm4yNZvY60CcAyoni4QW1jQ8rTmbP7aUANlujYSD7si0mN9cCBe6ymBZdOeyftkC5lbCkYs
N8GxIPcLEZFNe541bGyciUjMcoESaxo4q+qSidT0C0dOdtPg+rcOHDS/LU8YxIdRaCeZzes4nt9R
SJoLAtdMpTSxStgGAf/tKBxcU/FRqwvu1eo03fIyv1ZnpIfN0BltF6ZeGVvhCK69xDlckG2Vk0lp
cBXF4Ck/1O7Ww7enNrYLxYorgbSGZFwenzgwbT/4hqtXW5e5wpInSgVmWCb2f90D5FXMcEUYxKNS
AcZZQ9h5m/2qlexSKo64hwjNQ1M4zwMo5IgRMqRoyFWQo5sjGEouSnB8EaDhR/gpCgEkjkvrH453
erbfU81pH1UnVh0rSJl0vNkG33RdhObSexRmCN4atyXa76o/Z/D7OmHbattxBjlbPQKnT87VOHus
Waee9vZqXnX3XfrfzRV5ABXrQDzsdf4Vu+P2u6LlPNV2OlhK7TrgJ+KuqrOzDP4BK4elDL2EVJ3W
ajnflEZEquwrh6Ox0pfc5FaMv8z9RbGj9OpQn4zoNDfpJyzTsilqGotdaVBvY8GazZDh8g586EfS
G6Iup6V/7oJwZktekL1aTDZXsOo3LRRU1CNlh74M+WrdK1ECVVVC+OJPqqoX6qiNhLT6Y3cYlhUd
TlYpudvcys8I3R3sO2tiE44xDlw9V60Ihdr8CxApLo/lh32f+KWLdTTEFbwHH3xKu8HrvXOSa4pZ
9qFRV9DZ6fAf8mS6cG0jVBRnc0xvLcGSDPfR6ldZNyUD6eFF2ou4yDrUHnn90jU/rIIBhPfa9Z/P
bOxcl9tIV9vQ1ZrxObX3+36dBBJdc4YaEPQRzjBdTTdtHNwhPgyci+rXUuM6sITSsFTFVeDvJwcJ
fHcZ5CQ4adfeN+mJFqMl6dL8R30HaviAdOQsRXIab9xwrbMGyIbw17XQ24EQTLpuzZKIex3BJh++
qzBCIHOXDYFAZlqP9+TOHDFMF5+hjYN3K5Obw6+uiAiahmCweTtynKSKwwyuf7ya+3BkKIv4UAQY
SI8TJe+/PnNra+nwbIodxeBT3FtImuWBpqXtQMRvTLqq60T2oehmVO44duukGO3ClQkB7slyEAbz
dFPkGZ3M7fpKLAISCBnAdNA4xENu6c6mkm8o3oNdr15zrAvjuKf5de57UK56/HVbVguWLv9HDPbd
jKIEkOPBZ6mu0szmv5aoTBxC5j4efo0Cu54PaK9F4nBjqcqb0BYu5JWm3MVA+nEDc5UmVZuT5H50
wUcdFU6AG7EL8c6lBDCnheuQe4NA3hoqnaDHYtP98hjihJlSuphzzErX1r7K/IardT8M0ugGbclF
fvLRZqWqNq7nbo6GWqhno6MYDa1qkNEoc3X4t3o+Dt1lYcmhWwnXesTSI42mrn3rdyKGFZgKHX2f
BUQWqAbKQUNi+lmj6QWh5UmAxOfLc3ZZwS5bpeZDICt3HwtMJr2ZDOlDYSvcWHzsL2TelxS3j2C+
j87ZgdQx7YcWSuDYDX7VHHmDfe1inaFTQkwEf+DZMPKkIt4uN47Bw6gfYQZYKgyM+XnBmTINek76
WDlOU1cq2lDFO3kETu7CBYMLVclp4kq7LNocKm9nOkzvoOCuEI8zLXyjU0xgO2xX2wqia5SjIYF8
Rz6G4yNkMDNm1KNOVtuUP4LW4srVzhcCunjV8SrzOPwFeGATUZBYaUH8/SwURUUCY+NBalQ4hl44
0BZiqLga0P4C7fwA+iHhFI2x+DEvJLt61O25xC5Yr3V9LglBY95l2i37Edvqk4QA12mR3+J4buCQ
RHBH79qHuN0uf1AZqBiUOJ6PO4KHXUpXHg5C144nSA8DZzKbDDKhdh2jAnlVEj2Jx0gss4a50NqZ
05bFuQM1Ig9NfvlpJ9lqgsI7j72oACULDbGL7Fo4fK5V/xkwWjW9SumbM/OWuFCK6DzSC5XPDspm
jxNgojFTk0YdUasv2ZeU+DjeOp6j6gjlIB5ZMEzBy43Oet/0u75+N1j5bH7KHv/Rh7CyShc2V0Gn
z5xPg0L9gEYxQL0V91nbcVeXCuMiRzQEiikc3cYu2aq1/mwcole7RTM+PqhCFHxgPDmDXt2Ob8of
3bwmjoncSpTRC+733Zt4zZT4eWbb5I0KWfdSnUbtcS/0a6sZXiAXCXWZERD35MXPTqw5DU9sYOkl
CxJsAZNIzWomBaelIKISaSxMLNThuYe3Fg115tE+T9xEoXnhjpYwI3NT+2zVz8s1FudamrGiRkar
35bTvOYU//JXKguOgF6FiZ24/TeibNGTTmqZ8n4JR0PK3UUFTP+6O4oERciVfGr3aVsxU1eVv75l
1Bb8x84z0ft6QeGj0gZGswfgIM0Dhm3jwF8J8rmz/5/9upEtePVekn5J6bjAPqsDlI5PXrSZLf35
KUikS5t3O+ETrcETUMKwI0BqWkr0lW536Dftw+i9XjDDYSLLGjihCPGLV56TlYhG+IuSRe7sxFKn
DL+FNSxFawavEYavEQN/T6GIl+koCWYJ4t23oiJPfSs5B01vOuV6sqsrvMAzS0iaEmaqcVsJOyg1
HaXy4oNhHD9yPvaFDdzkcAH1DnSjkxntJiaJW2RzGWqcxeVdd1RyBJdGwlT+suUIgpId2H7TN+fk
PMiLQAoyQun0U4EKo5Bnz3MXGYYaaaSoEBscf8oTdj6hhSEDFdWBmVGXjK/PPEe62+sbf5/cQ5Xh
Uy+Yg0rw3oleGyW4ZFpBvVrBPbwLWErTzVkfJD2RjiTdcOcb4t+i5v3iu8VSO98agNtOI45O/1Aj
+kvLGtGSn1wLX2ihrjW9trj1b7r87DlTpUKbOJBSEfT9buZMzWcO7cZWtu915VuVrLnETqYSJH25
/C9b153g1lAOaf6TtqgzdRtRsc6iZtbxMpejm5JCRqHmNH7t5Q1l8KvrquUGEtkx29WNPd4RlZXf
6F4F3uXMsbPFruaZ44DahbK/OHllP2XCSavdkGZDej2gSNl3h73o1om9LB0li3ICTQwYw1pcV4JP
/jKBW7P3qlPiyfq2bb8kAvVbUmUsBlUrtuuegEijB7h6WJ7jjaaLpbeyyJFFLu388zlkqtmah4N1
Or5mB6wFndXnC4jDDpaw+wGA2aKWVuMnQJ92W5dLmoRAodiKcA1uF4qJFF/EMm7m5Q9Q0yGLLCrB
T+IULEtV1JeygN7KKcHAuFb/XB/i/kPd3LPPWepy4kPcogHBTSLbyPtT7R502+mx7fyEAeFEUpVM
8wtLzsmO4lbBSw29pOCUd+zCamdMrs+aLWnpKOKVEv+TQsgVv7s7UYjCnjak6bGdDqXZLcWSuecS
vlNlD1g49s+k5jsQvfSYTIoCmckc//aTz2sXlJkfl7+NNASjpxQNlPtqe8rSUQhiHmLt89g1GrXG
3RmR5uwrLcZ3oocKqawS5PI4FhSp+t275FUM63CeBUmwR8+cWVKT8i0p5JuwxA3zkDC177HM/JOA
9FdRhjvbA2gu+pfdc+ZFJfWD3Ir+bCCTZRla4co3mhh9ScUYbSJQ2xjDP3w3P/R9Dko8tXv05FrW
8+PVcopYbg5ChasEMHdIBX2paeGF5caugrqh4/ufSl4FRc3v+tgkqnvEjfCP83Bgouizj0WUDr+V
7RQjl91YxKasAgESSeYuTrOQyd7HB/LXIgHlshdOh7ILm99YIwtPJXrh2R5KELTvGdC0cGjNMMas
CzpawiQu60nb/7/zo8LsmmQp79kbH9wHkL6VUmLBinc4tVviNqCvDnSsjIyVGS/gCVFRIW0uj5sE
r9/80o5NYk0sIU1gJGbQBzeV7I3jEa2pAlqXqrVmlntUJ8Nb9BkeYKQ0Kk3L2zp0qMMEBPFd0QgR
uj/NTgp91IFBkz6xkZe76FMXf2cDH5SVX/r/jHbsMWQuB9NcxI963Ew3UP1KNr5imaj15ORr0E4s
P+cN+M94eh68p0GgneF6ja6pDayVZmQ2pcVtD6PC7f+qIMnq9Hvpoj4OthvUtIcRMwQc+QbSzWFn
bYdAvsSrmKPOaGtiSsGjLhuVem2r5VQKx9kvt3j/5Em1VcshJEP56Qv4AvCve7EUWysy+jzZNB4S
+q44YagMWoOTH0NjuZZ7upYJ8ragyu/KO/kUc18SwFKLhyK7xzPWdUBVTDYzwvKe1U644bqf3uDe
LjNzCntSeViIW0k4Q/l5QSYvs+l6bjj+LeM/6EGGSs1N5QX1tjGQwaNE7JDHohHCfErK800OOg+x
dIiy0CDF+H1kkhutGTAANYeFddSczfW4bfG+Pst90pBxxIn8uPVt0gvMCuOLddo3BPvR6xKA+QwD
nltNiDFgqmshO0GIzYmFaMG9NLn3V9S5b1+dpC2xmSBLeWgi4AoEMGExwuZmiQSCRarGjekoDiLg
7oyNWtz071TsACJwgL/o3t/+SDlZgDHxFvhEuFbsI+Nh0h2HFrACDniJN9/m4IMHf0eAV0mrkkZf
NVj6Lsl/750k34pJ9mhdL0FdPaWFHhzCsHYgxMZa7cHzwGKBBB/FWs8aRxYTv5nSCeA3PWP1FkZN
3Iqm202nzp9HkTigaTGPMLK4DJxsc8varC+EYdroVvb5zwlGuDMk8bPa3XnX0kNt7934M7JLl2Eu
QBmMwNs1tZVmGRjm64C7zxYu8fF3oD6ajBWSXVj0PNJOyu9LragMNH+8ZyaMkRw9K1isBtqk+cQJ
+TE6hoKix7zAsz5Ztjw8wfET2bDYPoOkgW4TELdCK8Pt+j7R15v9bMz0REAT8eT3XO9fHQTgPGEh
5QDpQmfVzPbsVYOslEl2R/x0ag7NafxlVRZttA4OXa3c4TSXodPKJYvdWQKlibl5fezvJdpey8ER
Kg+0w+V5tgIiU727q8bv6jnklwgbQ25F14xR1m16qSob1hlUhzbKJIZcD1vveILYizVRcOEgrILa
D1xgV2hmRs1e0QvAlrC9pY4mPovNIwC+W61lfgBWf7VghCAvMTqdhG+mc666Jv4BGEiq4QKyVfnu
RBuc8EKGnlOWM5K8q79mjT/jNZx3JJnRq1O1ZtgWMOnLL9i9MVKRAjmk92Ngz6vhWpS+pLUQp/rw
ncQKKELX93+I5yQc0QHDVpshgb5Wbcz1JrhUJ6hw/sHZPnRp8JvNGZxpHgWxcZt2T4o3aHyhOyDo
b7oS4aRKtpgkM2gtfbmgVpb9Fp8FtP9hnFrD/in66FrlQd5Jelmb9ekyCxjaQtpGXnPnwqiEq+GH
jPdYmWPoZZ6HinhMf5a7sgJHI9+VSMxtToRzIuPZIJaEcZlrGozNi/tthrHAOmtOft9n8HGjr6OU
2CIQocvKeXBzh5C6LbEGYfoMd5uflpQd3sCcAg6qKttwCGMIc5p5+Qcrjkr1y7yZft18+dyicpNs
2Nn6pyhBrFyqCVaSt2nfzNCQayfHE1jTVmIuU5QMegwTenZOxdQPErn3mj+X923xOZs2QYL3M5E+
4iFswhsypC3bZfPeNUmhCraYg/QsJNXJyRohidVgDsPk0tG60DewqFjq/t1Mo3JQ5yRWf4/EjwFi
p+GRVFzaaZH1z7qH1iHhrhOrDbnTbcTAA/Q9qtX0TapCAvoNXbuPULgyDjd7SMzmxPy4oXkuRAJQ
EZ7DeHgVyG0ocaWqVR8np5JHwkxGwcVRomncz37ETLVz7T7t6fMqQRCpriLGiwXC3s7vYNCsvOeo
6f6sq07mJ2reEzzr4ZhlExkQNnJKniaDgcI4UupnMaK8JBiHbDC+8G1NC+qRQ26wvRseyRyFr2gG
ij1hc0nmmYU+FcigLDQSDiOEg8f64KBhzWUqoHRnH0ekEPeGGJt3i4Ul0jTNMT98TzcssrzXM+Kx
eAvX+CJyKGKhZO3clNSWW/r9FFbpW7j/iDsMJOMNGg/QLQ8GUcVXwlhud2z9xPOtidnC6CjQviIc
IvML1DGWdES+J1TV9+fSZzr3UXbGKq2hfWtYAw1Jb71YMWZnzofIsjvfrNXyuNkOI0oFUF1ZSQaj
281AE07K2PvGLCzvyl824vXY5eLoTX6fqcnO5AnQhVE9N1RnwrmCHJ57MHYXY095Gel7Nr4jTjhd
+9ZtCyVcE8Gl5AwYJddFnyogjg3JNTbLZ4oCOjnS7OxaDHQ3u922sVnufQ9W2jQhdAu0N/UL41Ug
OYd8ocPkfKQYM0hpDY0dGrKa+3l7yHG2zJwKyQqagScSk2r+z2XS4a10RDfz+dFxzTEHxAdiembO
vZoecb4ek8kxvXv/pK37D0hD0Sg5Xn8Nw94VJshlNQ5vGYDdV/rp1M4L+AEFe5V4Z3IpbYETRU2J
LgD73TwQ7AXCQMgafHs+3780XghiwClBdqeEypBg9IKo2tMGzyzdNw+OhXJwgwMWSoYMwM9Xy5f3
IP1ujTACbtvV9AVGnzcjHs1gnXFwIM4kJIDu4SwxY7UZBZr5BvZApzPPIHY2d5FjyE+i+GYCFKg+
jDLF3wHhvlowxTCEgBKTpnkDnoegoRf79DzEr7INTJnUa8C3qyittxbLkUH8jXJ1ZmE2CM2FKDGi
8Y+904CqHU0GLPmIiMDGPpvXYu1MF/0Hx66YsKoMI4VXhIMaEcFTJ2THXh+GSarJkDhkGKYF/i/F
fanNmOIxcViyghQ1yowG8fATfmDernXaaUYSuitXHI6BwqCmRV5BRiEMtnQ2YKk5EYoy0Z2j6yC8
wZKeZHrNMw65wBoVDjZCa9KIl/+gW3Jxc36Uaw2PltoQQfwp6nwUHqEtWkV/4TTAX3OkN9IjT4/l
cLWFCwa5PMF+vbsCQB/Dho+15Q2B7uMxVseRF2dpJns//o+9u86BI5i0+ZUYdqoCGVXicd4+D9Hb
ZKL4OkVoH+9t4VK8num/G848UMsZ6Ylo2tWCwmSnz5q/6DjlXhWaCUA+IoIm40VXt2DMNnokDEv2
E0AYT/+IFH4d+ld5H8/tcMQbN2wyhRdF70Hj1AkG3wdJhBYivBMlgsphAe3D5IUmLQQ5l2LTW2BJ
SQ937ZyYArALvfgJelC2wnAay9Vt7IHYmvw3rnpHWh6X583oHxixed/FDyakx2ZurE8p4u7/H0p5
O1Au1QOjg7Oa5SoiKI4j8wqGzHmI59S6rgUD/tpoqRThg9mmOq7dpapUOIamgkwsGvjPhn1bXqWE
NsPRWEg8D/cQ0MwiZTbe7QfGup6kLaJ+pBT9A8CFBqCOpcStmocLe0g4k5F2JNXht5Rdcl9ZPNK2
qpyGwKdRFx+qpo7IsdAsh98tsuhYtKrfA9wnjbjdFduXdin+hPvhdywe+5GqP40iyHVnPcdJ3duH
DGH7txXup6AyCsLrgSjUb5bq8gIso6AtNVSSgSIB8+8EGbPe2bQGeM+ghYk65ZaWQegJ3qWi34an
6Y6LLpTfhzm/sd3ONs9NjarzRQLglNx4hKIIjqfvltQNmvBcljB95qizWbHE5Oh5YyXyxDXV0LnM
oyDXxhENmC1N2HmFI+HhpaPjb1Nq/ezgpGQHX5oLB6RFSHXnoh2kKT1EvIuY1iF4BRNWz1mCpa7b
WTcnhswozMEYEinblRmQKvYc5bC7dqVz/fF8EeYz7EE+TEbcFavxRmiXZlolK00lwCVDz9gbholE
R978HNy4Z7ntNToBQKAkVyO4fvY2b49pO22nHShJk+uArQjOXWxTzATK8UHdBksFqs03OH5iACAM
sJ/R6GahlmmavEUwdp4NrjPMWzr9fkfGcJvMae1RJRUTtBou6zJ/P7PctAxfE/inxPAOh598lsNt
4s2WAlRJw8tFsK82t2GyoaO/c5E1E9uqusNhCCQwpq/U1hYTvTAkRhta0oEl31TXvNhh7ZjpGmcu
pd9zELdprpsbqkDyoPEs0RuLspktO/t9sMkT4E/PMMvNlmpJsWMQlLhEH538THQLDIS4nTDcdeOK
x9vTcX+NKRNs5YCwgXnQXYBWRW7Q4nbIEemzhsepMoszg+hr4bB6i5pobw3qVBNGN2CYgjjGNzMO
7yv0P5VjpUyW1RxcH7u5qmDMs/r5LdGh12wGwdiD6Bm3cfO11YrhXEu7rzAdUPQt27Zger5H5+uf
cmoYjt6OKEI1qN0ZWldegpdAP4oYvq8Fz3jOLnEPDskXhIUsfH23YrM5Wt/pzYbtrecZNBM5hXBW
fQtqZoNStZwR/1BGZkJ2n2CUGeUEFmqf1iX+kalQ+KJS+lFRTyO2JwIR4lH8i9L9QAV/Ffdd/LGU
J/QJsGHyxXQk8DlJzG4EsYvXpn7qDjVkuMBGT7/JLKfg7j5Y8pScgXwNxW4EuqbgSN2asVlUvMQm
QCesu8H2cfcvZYACoB4KaUfkjRzBwP26KNsueAO/pWrDJ2Zdp5+gVLO/4akU2foCYNHKZDKjnmGB
OdwT3gQ6+dqkeV5Y6e0FRoPjRvxa2nPIKz5eLlnftd/4vyVGrdqRlukL4IfDN22u8tjrngWA8yUF
syBRb9980xiIM6HylGBUq0ueSBRDb+EhjgiH8NelsO8UbBZ5SDMHZ3/NMQm37maaUwCk1O/3FZre
El1z2yWkgvZz4zWoUbwoUEuR4AgWMgjKjo/hh4qbaYC9c4q8QTIB+01n6QZSquHo2CZ1XDmksu8q
u8pVBX1oNw3uqxp7eL6yDa4LoK4Kzpn9d8DY0GbkX4n+aPwLEqeqgNm0WEpPQyYfXNlp8p0v8JTu
4nsk+c15JxBsFhdd/KOwJ1YGv/dRo6yRFHZO1sxLXtXXXQh+Gbv2RKbHjS1hG1T+9TPzXT/50lWT
NA40wUrZvy2nw9gNoxlVCU1VQmQ6vDQ3y+BfSmAGmSGIjneH3SLVg/y5B85vc5xEaomBBuxWiEuo
jCbTy4FKPw43IGjRwzZGuS4bxsThEHp9v0aktOKZ12ewpSdqHZXF5y8YKTNP/CsWIJbLFb8KKegM
J/879frYqvWlb20X91n6N2aHU4n4jCLjc116IxM5qbIJGEiMjocLrKWU+Zu0ExxNLoSoa8lwulOY
5J5SwIEMUruRKTooN/DqRcDpoaHDT8MM8Ke8dBmnzhwx60WE1eAJRfOpGXLP8PIESoEls0NeyeQ2
Io9nLNJuD/BQbAKzLuh9mf6czxtBBRJar8RQs4uVLuc+aGon+WNHwEY+0FE4nAkyn4SFpvk2Qqke
aVzVscLDusKnOFJmIiBPwtuEklPhF6Rk+G/HdRC0vJxbXJQsXrgQ2OlzMNWpM6Yjz9hy6TNnwkOW
Md2Yc+FRJjcpBNQh4tCPBmzZLnLjrYZlYceBMNRKMikLZPGiG3Xt9GrXdBDiUHqigSmD/4uD4317
MOqEX9r9zc6IiW7kOQUm0qflXzM6+pgqBaS4sS8hvgnOTyYq5bpn+Cx8WsIHx1xuk/xuBLWzxInr
fD91B+Q2wAE4tQQw9mk5K+gwwxLqIOeSKyHoCeZJDdhA7QYa2d8UzH3xJQOHZ6XYx9cU9E/4OQrD
cORZY4TUGaOo9ihRVdTcD+6FrHwReW0ymo3crUWBtCZGb5dG9pMdAxJd6NGMW9q5kEiTb1SkX6fH
DOg5Om+Oi5tHMDe3eMm3LW1NlfaYY32uKHIjAZIKuqP1HGGZaATAv13kelehbu0OjtmYLZIbiE3K
xJp6IeecypsjcvO4HpsOjStWHuU8y0dE9EB0LAdeUuSDF0iPTHMleoo2fzE3oMcx3gdwtMhq4D1F
hmZR/azvwbWZnRbVnNbowR2pS8NRxYEkpCEzz2IhiV9gtz9j9zp4s+OSReQhRU8cllYOW1gwQjKD
PBrWjqF4TUbG3NbMzC0a9oCbLSkITpA93vUGoojl+co0dgOgAGQUcaNqYUSXHFm/j29ErCdH8FM+
OmNOk02yHgNd7jrZJjgs/GoWE7PmOS4jkvumkmm0vQ9E7HaCDRaRiZwmeIETLHbOM7rjXLavdKcq
fFhf18ToHGTHd0G/LvOHLdnJC4dWt4mmHO7inRec9I4W48HhhH84XnvefG0/P7/eYw4tIlKyYQu3
bHyHI8/TOkijucnAcCjZ7p+tmqMc3jJEdKUHh0fivEeQ6AtxyKZKhvQY0B+SNX8ZIfdQbIGUcYh5
MT78hB7k9+RlTSOQ5ooixEwc0bk+w/aDUohoR3ETh7HFARLm76tsHZnveAm2Ulzh0y7x1yND7CdN
iA3X0CNTl160jUQFImEmOh76qJpZHLTRQc/NE2uoA6HVXqb8s8OZEvy2SsrBbM9VSYOtUyXXg6cj
I+ipGwaSXHoc/fCmwwC52uzMMXA8+E31an8KvMFqX3c551zj/YIo2Q0UY51/kGqFH6eKGOo/YssM
Gr+8rdQWS8pzcLK4XCAt1GKP8HD91gD32MOrh0J1pP3+N67hirxxEHcIv6ljdHv/4DHl2mpQtskU
RdS9RxejagD58cXD2+R/YO8hrR6dmkEXeQ6Y8zmG6s4izByjEmiSJnazqhPlTPStylW8MvYEkYui
JreY9j2FNObfxp271RzMZ89suWuCGmn2ZSOURgIJdJiIVq8uDUT2xNC3KxvQjBYzG6OW3eqU70+L
gDmaW6U8gy+IukDZ5SOtvE49FoU5gkpVbpFHXsMd457RRxC8w+gKAcj/cweqh9b16+V5PJkUtfAu
D8OYkSh1Fpu19R1eJYxjb6+EWu3LWiYXMXffjAS7pmmlk/NiTqdmea8YXTL3OfKB5/H7ZGnrjNQk
BX9DIxuW9emirQ+xOSBRdefMbY1ytkaI3/Of1+si0hxwC6lJUGqfTVKMn3iUfzrnR787U3A4L5HO
AGDm0iI6RXMxzhYnDeZH3sdXzXSn/RlRNAxN+XLNvXvuItzUpRJyhXlrjJV2yif4NUqHYS9hkcGD
nWwwa1EwSXLtvF5YYUlXhkQCMBZyXK+TIf/3bgTyAQFcJlchEJnutQahsrW99XYJ8/DXkR3C8W1n
jUWjWJ0xXIVbjRnja12KuRfoUuEdx7yL2atNDpOuH4Vfw0S3L1zuzCvYdXjV2LAps0BKLwgDxB8R
ICchSn2W+9TCZx1zhG/tVOZutg8rmmtzE3jJtB5GJLajHXILavWBAdUCq1eZ9j9fyARoRBtbS4D7
u14w9g6mhPn+ZCBcDf36Qpz9vznVcDsXwgnF2mFwYW7wRwJF9rLvFPXbr/GDCmLDQQ8HCEy6wlJe
ZLRrbR7v6POH+V7UongR6rS3X3UfoLlAghHvfPZHlFEhtO1HUZqnVBpBMliutRJ8DdpvDqIXwQWt
ic07U3uJFMtgj8fqJciQQsFxxQJXBKH6j5RDHgFI3We3M+dUv++rTgzaeFBjpL14qKH92kLpKOOx
uX1YXBajZQNGSo+r4qOFfyboBgHZIo8MhLgh8A/ktoUWQqX5XUymyPSO8lQlIGSyWy3wHFu3ejP7
yvIR0jtK2AtOpj05I4LVAJ2fIx2gWnRPA6MZxUULSTKW8UCEkcnDS3dM7dkEVqa9OYZFZu4la+eI
hShmTguA9a2TRznrnCVypmUxH944BKO0UT6lWE9CdOblHaIICrL89rrwynuQzr+M89Jw2XiMv+Ra
Xm+Gx0SBXmdY197AqLxQJCk6sXKk+9A5qn63pchGYAWp7ZTZ+nUADbZBKcKC8KFEf2f6o4n45VUQ
/Ys0ydbyIF1JLpERp8hzorkW3DfNukQPplPUYurrbYvvBbSPCkMYAjhAATr4+50YNsF0bZurBjS7
tdL8oVp6eX2p+7Iq0x5omdDpOJqlgKq1FBSFJAMoOlLawi03Z89I2iOWGPQbdnSE9DiwW/8pBBHD
c2mHJznScW9RaAkVAGNDAuC2V8AqE6w65iDg+c21h+ePh1ZsZ0v3CxGi27+miseT6GQAg0PO4fRJ
dyt+sNbazhWZT0IYJCHuttpOYZAAeDx8toDbOOmynzq2rupjT0/RPESRRoAyZUNal9Oz8UC2tKji
uGF3pxkbMjNQwFIuRYd5dsQir6HoEQRql6/et0wYlTdjvqVTzzqc/2jQa9anWslgeEHNXKLMp/w0
Xg1E/BesK7qQCILj1YXBQJFfvlqa78NzBkqGJQ2iFrq0uSktgLo8Q+vih39DQtH/pdoYzvRaPOli
UgDJAe3brm8jEB7RdbJGge/TsSluFjnJ/WGkZ9cjYngIn8ZxMDriALS3Lvrq2Fne2pLWwjsLG2mC
qBB6hFREHxYMdVG0wLN3jZM9mKo97I8lWDz+8L6Fm0uJq34K1XQPsAlvYWctQMSWBpHVhAfTO06X
/dquKYeFAZzH2qg3eAnUjffTRgGLG0k2lJNnkqnExlPv9abs+rSf/NXBKVzbMdWSY2GSikwuTkCO
t6c4bhzk49pNYkwwIMPcXhjygQ0xz6bfCh0ebQzCGK5UegEdbgS/vL5QOQ3t91T9DVXOQQ93lm75
p2+Wmd6NufX809nwaJ5n7oW1wpg/2grFAcGptCEFDt3Fz28kSCr0X4yO9d7rsac00Gym9LMe8T+u
kJmSoGD41bsxvCsa0jshmWKWbJxSHU4RVGdzLkhPH0Yem1+x9Xs7lDRMA5+1jMCqewr7+P1ZCEYR
14CR5Yr8EqqFDIW0oXR2hR1GNKWObPkk86Fyh6jXZBI4p5zBou1/DgNldAJZmpYn+d1gJRkFeGKZ
Z0WIrLBca8aZZm7f5Z1abaw1LMvyr9HSOsoI2DfPKCCD6NZxjWuoM6a3p1UfVU6NqFVrcDoEynf2
UqIaVM2rq9GfKRUDcEBdkVE96RJBmLgSFrtTwhs2zEZWarhXluipL+s8yGTxE+ZnehjFD8Drh3Qf
4z99g02T8KM0AnvvAeDq5oeUHXsdhS7zAccRb74z7rBToBzogvqioG3i31lbfiKEZabLO8kQsXOK
PloEFvBFqKg+cHPu6uHx19I2t/yl+iXvtQqEV0dCJOlMm/qD1zqvOeDyTJ3t/kPDHVbA3SYoDhhT
8kE83/iKIrcfdWTzRX0LMamz50gKwzRjPKm0NM3VXfpkqbLCKyrxtOpJtam40QI/ApPzDs7xSlR9
McLOl+bipTV0j5vYTFE80DdsSVJXC09V4EYnTkkY83Ok0jggUUfbMVq4qd3u7aQg9pgjPE4ciwrP
u+wi5PmqPx7HZrj7XgJ/GAkLGu10Or889Lv6BiefeqBkf5jCfjqaJ4pi0e/pzVhmEwLvP6ST6Tub
66xCtEJA4hG+MdF3pcYs2iQ2Zs+BYAd6hf7iCUIJ9n53yE9paVf2yanqoTuQyt+3HY+O4KfMAcfs
iTrneXaNRz03Au1oPS5gA0YyDvasv5vyLRhyCjy6cSCLGukgAwiSMkBicPlD2/QXmlnrxJxaPmM1
SZ4a0PH/+0J9GXWY816mYHqcBtaWsQubWKGPWDoQtrssL6wTxwLHTYcFr/17wjLrxdQduluxoutI
utxo1QKBJ1S8vDsPORSvDDLUtc+zutf2EwNcgtf8P70crRoKVczRmSxqF5VvobBbNwf3p2OTYCjJ
0vqPQNUmT/VmsFekzDoEWaCBp6xsXGkQnueODzjPXxiHMn9dYip6WiuyCM5iJmqRNMJ6jn5YjTf+
FjCM+FSMuX/LVAhAVUV7gfqkT67WfEMHPNWZ85Jz+pJes5PDC5M3pkna+dWbNW9Bd0LaYUh+2Za8
aA5PzfDk/qoM4gaH8NjWyub7WkAkbHe897ghjg3Kw9HU73fbRcPB478kCVfQHzoqgMn1PWMeVr26
r2ecbr4Jy0x4KrNPJG8cobkIStd1joZL0IxIMszJc8zSP/KEVIPq5KVc1t7J1ryNr2eqERsQKQJi
7SsUc1UGUVQR7PTCCXjpqJUnsq2DqsHJ/x5P/0xG2ML27VHzrEUXLmd2F/udQoYBd4NCcQ9VXd9W
etEx1rgrdDaaX4qYs5DL8cfTq5252MoArj6VGCDTKz2aOrfcxDa7c05ZR+V6Fk3T8eYpl9VRZ6PY
4GmtlLgazKZ2EXRuoa961YLG6+94iNXW2vLANjCqSS+c33WAqMDBQUE/yvIJu0fK3cHsVOKWh1h2
11CQOSnmq9ZsOWzJrp3XyeJYHXmLasd9e0RIYWJV/xipRcG23dgxtioIKFPndgs+Kb4KS8tkoN5y
mDnRYMbpR7spj/9TOaOt/NaUPGNz2D8X1lfKY8cxwdB4mn/86N2C12MJdFR4T+I811b1h7Yk9jF/
dZGj9/lfOdhmkbDoPhrCCCD8/AlZl0v+gqchwTxLyl6Ks4MRDvbEoSX0/o+mf1ktk4MF0nIkA5qH
Ri87oxH2cxXt6YaX7ZwKVCHIevqAKuHCYwJQr4coHfdwTj6y7XLe2KVdUsQWPVfl/7kmLIFnmXVm
RQmG2rVMFHNuqANPMmt4bTBESVkalkq62odtVfeanuGa82oBMDvCs1w0vUKoDRNvfrVmKOga2aKR
yskho9p8s5IHeipv9nlQuHl9kLrmycHudgiY1DYrIQnGprHwZnt4PMbSI9c2b6wUEYQKo+Et6698
QHBHPsszSf0KJ2g6O9Juabnk3LQ2bSEI7M52qbSgMj37fHy5VgeBEx46MMYrt49ukXIeuxt79wQ3
47fnqgOdii553nEX70CmRZv/IrabBb5bRvOntfrqyfpyluJW8MN3Klkc6blinafx58H7Qcv0G7bF
BFmsdEdujgKS4f/MtTFvrjSNEBqSe9QMc1sZua9EUf7Hdsvc/vELIeWoxeHVxWTOfJb6yFseowrn
Zw+3LpaOsy9wo4zSntvhOwDqtfcWdHjCGJj0m9fbB+/MHtKNNr37gqiFxt6fVaz+3GQ49O9evU9w
GnjO/BZjPyED+Z2QSb8LOKOBxIpFIISx8WCDXLxaq0NeTOfwTjYwQNJkVroJRs+2nvjrPtanwLPJ
FvApXFmGPTN9aIpG+g2LwqSHKd8KDZMa5dt6Z/NR8RFwtkUnoXz6Ihhdkicow0vJh3RTdwomUTmf
ybqBU2jQh9OjAcRy3Hn1tIpvkJfVNHd01CZCWEI2WLWmUw0mMcNWtbI793foiXoJCTt+GT/ewSSW
BFbps5MZcSqACAvnE6QRflhIG708oqMlBr4J6YbmGi77GhMgq9oVN+/QJXdCdMNl8Fo50SmMDqS1
yjt+P8wsV+NhjL03Ecx709EIuWwZxqiHpwWC6HtS2ZF0MveuMiHClXv8CveRmbXuNyEk5xqkx/dO
S4iICTQKzL1+kjjfYTyxzEldZ0vTthFEwCylucs2t2yIMEh7i1JYLRCh7YrkMQz2Qow7y28fkbwd
qLYvDRvTBBTY/zyA0CxxhlZ1oRc8UlIjBRnUHeCwVlskPpzBpTOitG7cmR15hUTnvn8tof8Rh/yN
SGGSG9nFnztO/I4wozjkbUAXhg08TwWhM5I96KXnaJGBWs5K6rAtSXidprAoQDgZ65ckz+JusBVr
/6dzpN6J0XKUM7zkcAu56bp0T3tZJbao7KcQ/qCFmJZ3UTLFvqUUCMd6TL9jSqmpsu0SYFuqLzTA
oM3KvpBslYWe3SJiz4XefmRgc9eYVJxGE2o8s8TX+Z/IhXE1Zsps4QSpjFFCoh8awrRuROTm4PHo
2nru7/T+WMPW/WM1GFr29yEo8zyqxMTCyoFkZpCXjrzRppiiCbFpGXfy7ATONY9DOs5tTefhKRNE
KmJ2luJTrag6/FoBPHRSQ3tpY+yMMe2WKtoAx3bYhDKcLutJxOy+tmlqXBMzxwWR+EIGxs51lvlQ
ZQ8926ldjJSPezXxY2xUKZtrJPyskMv/faTjPvfBtKfMEc4L/7+Zj599DsxYlu2gTcMC6feGpp3U
4I8lwEFpIQ3krVTTMNYWm1anB3mOC1hUPk2R35Yrco69xTYjs9tkdrC10v9kLS+oWzbfb89urzPJ
67+tZvNVhH/8V49uQ9iSjrn6SXSxqH9ahQvxvPnp3Zqh2J2Qoo79eVqjVySVZfB6tRla/OiKujis
kAYkQWrGUEsYvOSZ9ubGmbjHdR5PcArSvwgHPtJpKNTx2e/yMqtwktf0l2CUoHYczWHgSWnHxgzr
ve3E2Ey4o4SBNU765a1ohLkd0k7XzOhBIEmAcrl1eGLmdKpQq0uzznamtHszMKb1X+PLEaZlh23v
KHXpzzzrOcFRZ8HKe3UKP1SLVoy0rl2A8O4gQUD6EXdioUTXS/6BPRXcFIl465Pgz7nz4Ff/ADCU
NUYs0w9BwEFAFGnRkuifJ2dyY7a7d2SRWiuXl/AUg64PAZ8CoB/mbH5xRhABHEpAlGK1iLaPDfNf
OnlRglb7cRWu6VElpDvoCyNCJ4P4nzjySRCamMYb/V9SBSEnGHGwRmhJDTPPApDDEZQPeedu1v5P
7dmLw0gR/OEwI9LlGsLqtYB2Z3T0kh8dS+vvgDTOtlRv8ndrBwLyFwdckVrckRRqayrLMLzMtoLG
QNT/6UXaFS+9LPTH4Yf6p5/Eo3KZSQUUFBOTTUUHQHr1WsF0mYpcfrVkexqlxs1RiTQF0RsD+ams
EGZ2+5A7PD59ws6LdQpT+75x2Os9OTwPt8jQstGVIwhn8c4dSlPntqxONAayvwMCrRN3KCkQ/gOk
rEzcJVizH2d6A3Hr/Eh78y9q+936qKFmyKix2K890tWbI6dVE+rq5RJBfrhgkeOU/U6LJGZVrwjA
hx+4OHqVkGMp2p1sNqv8T8j1RJYsR49OOX42MQcUPse7rSWvbHctPyCWIozS3ajrVL83/f9RIIYL
pJzqJPqd0l0prKfb3qVfLrSOZ9l+HSVpIATmmIzSRIGjrv7k5xJZfJB7C9FKdUlYFINh6JLQTaNV
YFPIhq0okVqzTEDY8IGEuRs9if8gC2w2XohkZNgMEI4tr7fMsOqE5iRW20YN8KiT9mFOWY4kkxGE
1mBJ9nIz8cyuG7uWEqBFJ/vjJOtj0XAJ9iwa/UdOHfE/x9qtAZyQE2JEBhzSufugpKXm4SkuKuRd
jKl5OdD/LXg8rjeJW3ekirTDkw1JZ4/Z+8zX2Jz7wJWufLnaPeSabWAti22HQ5T2rIgBi9CzPLG3
yQCh6a3i5Qv30SmTl/opYWPcOBb0Yup2gtiRf/oVhoUiiEEhNvn1fFrLHuEeQ/FscK/ippNHEplz
RRuQq+Z/8RvARNFWFpaYmCZXm04XFLfVGFjkO7gvKRqaEuzcUY6CoYvxqfK2GRcgQoaiYC1z0d9t
9En9kiWPvTvqWve8xZAlKVYuREjqKUZn+tr0M6ySBt57j28bFEO0wWCxuMDJLrDYkJlLZhYmj6CQ
WBWP+kYcp1Tpniu59iioVRq+P4JC8qCrKSdCvnJs9YIqtG1+2sSFEkGUYyfciHAgHR4TcS5d8QD3
Jwd6H5aAJOCzac9xNxB+akcyC/c4luZPYOu9+BgtsZLTbDm3jwpAKSTXQG4+Ocq8JVosLV3HOtsA
wHRvdn3lrVKouHAJS+GMhj9gsHkBYOoZk7XXjMoQVtmJqqIZ+60BAaM3UB5MvX0yqtVk/ZT4+6fg
U+qDY5K7+hteT1NP1bIWVAA+SUb+Gb4y9e190OamQoVqA1t5e4miBbgwkB6fo+GcbjVCr0h5ORW3
bWlvKC+3wImc59WOyB8dXJLiJIuCU/ZoIxZ57ovW9/ne18TRWt83E57tU7nF4Spos6pIgNNxPB6i
Aycr1uBsTtJ+MiY1T2zdA+EuFjsqCtUte7he4pbmxicaedSfnD6SGEBeF29sO1acG13+jwFyJIqd
1ACpYtP5wfVshGsS/0MLgU9Bb63sFwIXxt9PwRWy/xGmclqLyxzK5yEYxBovXofVZVA4MxY4dKty
hXEzxVoOx5fVubFrKNN9mmBRq1jLvhTe3gcqsRIiULoI7bD5VB/roZ67XW1R39cZwyfvBEetUwie
qVw2Pw7r+8KrKpBkmQjxTt/YjiqjOtK+DR5walXDmChDzYyKuRAG/SApJrSl44iLxxXtXzU4YsYg
/Q9c6whK12ET7TEv75Aj6QSNV1rX0cMBoi6BIRKUIzBsmi9D6f66yRdMv7Vnz9r9KRtDDIxWh5n7
HUfvOPCjERQ8s/RjPtD6ss3Z6IqoyR3TBSg1wxBEhm+MZooqfwnB5g7unPLlqtgPJ25t65411YzA
a6OZaQC6hCI0HeZfuIxmBpAc3TVvB8FpRa77zIKVOxbn/imkKkT0R0p+XTiKn23cPYkIPAtjG2CC
I956vzWYFtKuV/sOnxCkgijHTCJXSmkD5UnptUQ3qn+fWGvkJi/nfS4Dtz6rCCCuLK+d9NT+ucPv
3wli0AAc2HnB6Tdc5AnJypbJphc157wdS6PZrAI3Jdxojwhv8X/BRgmwW1dSNhS/N9t+waDXddPW
TMGVFsrQLLbgq9FfKfyULtTmCUkPLs/R+jmzzbgcrz5ySA/W/k0gYQrqqefDqVu9+RS8fSUBJdzl
KwBTmwUMfCMda251Mn4eOUYEAnZFe44wjCqwe+258JfYw+BHs6UFfgoRPCchtf7OLlWzwW38AUYK
ABWFFqJs2nPcXtJYlsn6q9Q/yNxvB+k8qu4JYNKYNG82pM8BkXZIiBvPuMcGzi1yTXUPVIlTTLIZ
BeMoKMvLMEs4jkSkOuFSDw79kDRCAZBMmJm4Q5j43yzwlKkqvc7V67y54aRW+f99FYK47mdVU7Ni
WBmHgJdZC/DH+Zp8ytepxIh1oft4Guw8/IjyVurGhQGYB7OI9Tqnjg7EvlLEjiXvdrW2PToO8tS9
3q1dw5GtHVvEVS5NV2D70RXX7D1UbvnoXBkf5s40FzyI6ne6wVwRwNa4qor0FkutpX0qp0B5hZqq
BAA7gOnFhDfV2DmgUpO1adZ6QINsPfsfxbswlwJCik1/gf6u+4nJj3jmJ3SKXOckKQ5pZuIscZ+2
CUabRiv1gUhUNXkTfEuDOG/kgVYNQsnnGYp4pkZQzG24CwzGHQArBisajPqBDZTp5726J7mJdMy4
2S1SfmjaO1WpaMiMOO2lCF2SrNxjt3sD6pQXXiJcsuz8Py+iMsFkeAtx2bP8n3hJ+xqI05ujNXHt
pnLh5G0Gp85FsaP/+7bc0tAHWwmPLbJ9JMz1f78py5r24paFOdCa/BB9uwnoCWx6cz0EvBdYI51g
eLghF4LVmmjVHdaTKeylB6hVXwqn4whjde8OtFhYdqPLEZ6FqbRklfSSbMpsQi8LAurUszoY78Gs
c+WGQLiSq/BRmthl1/JL2KrbUw3h77h/LbXbNoiFocZKIKFyis2P7HkhsDiCRvoSqhLYelpoBY/k
outTslHu4ihyqS+TS3AefJioth/nsJg/xq0w0RsUOmhzWO8ki+Xi5dg3CG1I3OX3M9ayIaWnxknE
QzNFn/Hupz+scltO9RWZ79IFLe93vTVqKTKmJM+xlvUqLHQHD3PfyzL1VHa2cj2muN1ASdHPNM8g
Qc7vmcpFFdMKol9vNY7yyw2MMNiyKgfVvutlv07ktXNZleyD6G+7LDqvCRHBnQs+SndQwzqOlz07
fD4dLrrL66bGgIGHexFzwcwNhDX8U+jWosunZBXJ8uvEDYj7mbof8Qxgsy/HG1yNcucdv/3gO0ro
ZKDm05dJjAlCPcWVyDz2LMqPYexTwaYUQh5V3dt86dKlOdsPgfzshrKaMaozKdGr/7aga/z/+pjK
Dd6UZ6KiRnTVRVGqnNk28tAznYW9xHbqbVRCjKzfx0nudIWMHkWkWEGsg+puyvVLCqDmimEZBEqO
GYipR2mbwVf+YKui+yzhh1mNVq81M6kDQeg1yx4oqBeJIDYobflXxYkg24ESpoQsOxTyvvVt462A
2se1hBtJFKUdNEpV3V/ym8AuDuw91pyaXqj8xBN9LYe7Olgb64LqbuPPQ6f/8kZ7xSe6alA49yep
qCmKP9RlHCg+/T08i+YtZ8F2RneYskc/MOvDpVwmmkg44jiRvOSXE9dcQeB8Oi4Ach+n3FY4GGhN
edcsm3y27Dan41fgAfEoUttk5ekTIkd30+vhYYjgu1sinK472ulPwv5qnjRCz2gmp3VZh8ezb3ms
/fWGIOl4UbgAjC0DyAVzFCiC2TOacRBKv2Ho7Uc8BiWiJrABcf91FZXlRibQVUqX8TzUZOOffH2O
uQuMYYn/XJ17ju8Gth/4hxBiVyMWTWwC9Q23e6Xw6lnDJPKAAfbkORLoXd0tt3dIRoT8RKL/utRn
srV6LgQjuHE7M75Ka+oZu1TzKCBcnnkPWNThQ5+8I2FbaABBKCuQsnkibONLBunk1tN2z2dWtuFy
jD9kSs6YU6p3vX+F96Zd3Gu0ymQcsA1gp7QZgBtCDu0KAludUR7LxXjfjFsc7BKMMcIMFjcqoZ31
UbtbxgCUhNwJN/uTzDxHDGa3hF0liLUE4Pf0OFpTiPpqESGUirXIp+2YBHhFllJ6WHuo7xNrDAX6
czAx6qL/uPoJHu8eQz4dx7SVY/PPUNEKX+/D1Ra756eVbGCCSWE2/aE7zyjY3SeaUK5NGK5UkDeR
iDr95H3K9BnwxEKVNNzUkA4QAeEjHP0LeUy0ezBWvTAmUc355VnCugG8QlnssrhzDD18vJhrVfqO
dpAOapweCWY3jNmx+R5026taHpJJngl9JFBEdvk/xDTcNNg5glr73KugmVHxZePs9hNITZm4mUhU
f8xltUvoi8I41XYiJr+/uchngiW/w1gJ6KZJruzMCqY2r5yQsGv5qgE2/fGBdjdQQQnnKbIyEcpB
CicuRtiSr6Cr8bFYTJX1Pk8EvGRNy7JYJZo8kfab48j/fiUwQS47j9vEmXPVj8RxK+rBy4vhnS1+
FJHp88Ryd6tTTQbeUxjdyQnPZ95JnyP1krmSJhTZWKBI1jKLfNKGbJHdI8zahHY0MeIEDULSZoyF
vU9YVB2q1sxx5woYrk8g+1zi5m/GE2j7BdnNd+35waswF5/YMse0zIYJ7OvCqSUFCy1BK7gEJgJz
ajGd6H1a6x6DFRONjE2EzLum+1cnSZWOUW6xqLQdBAdbBasZGCSkosfwPoEKZcyUq9SVKqUtaTtI
KncjwPhLxkzbmhKzehicUVJw8BCBOozJj5DQTUaCM4qb9mC5ZafEmHHUUH+MkhlHrEeb3vAmMTvn
qOxFBNdszC3MLNh8+BkeHmRC0Z70ZjXX3K53gE2JaDrIjmCFwIFUe5Q5sh5j3RO3I+6UJmtodx+K
yXRgExWmRQxID4Nw0AGk6Ca9TDd5LtNf6bTlc1dgUtMb7Lf+o040ohTAp5/z8LTMf9niVLvfxV/u
eJr4zPjk6PqvGayMzmz+hXc4NowRz5Lv3lehxAUscHPjI1xCQg6o47Wuh2BVxKzzkpZrshzz9MbL
1mvU3BtxWivF/y0ImgS7It6eDXszdfVeKowZf2OwDd73Fa4No8q1kBC4FPJXG+1BopEJecruIcS2
56sJZzIJSGqyUUsllG0ILHDWiOIdwUueFgDV9pqNZa5K7t6R3xLlAD7KhmSusWwJYb+LT0L2ro4t
ucr5K5j2sp34jRVcmH9ZsSyoGt+z3AZiUAAYhyUzRhuYd38QU4T1KTTcp1HvP0rmBc01PgqKOPUU
K9fv4Rl3SnHRN2lVSXTw1j3QwTCirVTyVVxwpLJGSXpav2KiM4Jul4p8pKk1nC+B3HBo1qWSQbpk
MNTf4OFxp+jCk2i10Ee6Imov3NW47q85tku7Ion/NdFUrTR04GGv3zabpmaOLc2/oqQ4S4hQq63C
88D1bwIgiWiaqsv6+6rQRcDRdJBf/UQgMqIBPKpH9UZCB3Lwl+VouxNlWJz/WZ3PBVerLlmkBm4p
pKzZpfi/HwbD1WorXJx7y8pTWGJw82BkkM0rGjl2QIaQwhxeqkXT8iexBksAWP0DtOxfxe7MA9B5
lBaeF/MbAkOW3Z/B9irzfqJLjm12GUryLMdIzo+f+vp7TO+hlcNpqvOYaNHCvcuqrEVZ77mH4RxO
iL213jXEBVKlH8uB7OVrMGHgW4Qpl27iWrIfwL466kuHIiUf6K0Nn8B44tZgSbdAyVBB3i62/a/1
OPxaBgpKoHes/ZFxCd3d9HuVJJb9MNmndOEcDAUIe7Ak0XqbUZ5YcDGCJRujAcfYgUHb6oJjegt8
u9n/Weh6Tf7aETTUSIrFWyVGv2JBw2IIASFjHxRxdfhRII/8umHDQKFspMjEKphrIJOpP0jGPB5r
5TKV7PzqtJbwQZPYOkIUHXRxcZKM9dOdUKXwmP8UmaeiODypYLGIgwH+tSp/hw2Nsv9awN7hgt++
0mYJ/SW202GW1KsrGBxh9kaerbBXSQmQPFiCrs+ga8baJTiYqv1HaxswSgd51Mx3lh/yGHE3YBDu
5VPUBbJnRgJbFMyV9d4XLePDW60LvapW5QQMwR39lipFuWLWm43QNXSURumhx143K5jEDppYGL3G
QQen1E5w/euPATp/hjTx7bzfYCK+UWNIwlt8d/k8sZkImRcAVuDWBLEbAmd+Xg77J2wKPSapoWtd
zkj3Bj6H13Iicrfom//x3qs7Xi9qKjO5ky84EWhzlcgmyCCfSehpE+YPV+wTs0Ft1tpoY22dAM9a
oB3Pj+NkEntr1FovsCjuni2MLBRfRooarpL+sB0wx1AzaPl5RbfpYkEgAULVtQMUItRu/cMVsGkK
vhi6/s18smZeyoSqzpCZvzNxVr5y0uCXqU0vb2iVsZ93HBNga4ev2AKYqL3nKwFdf0pOfUCw+kqm
hXD9iSrJ0R/qooIWjeB8E18cCgTHTIvw3ym0YYi6kMQC0mMhLf//HlLn5+9rMDSvK6mzqAKFYW1U
k5k4MdZjSgSy3CcSYHK6Lj0BDw3J5kr8f2qSzOgVee0r0d33SzomJLxP2ISnjxUrPO01h+K+meWE
WSyIufUvsFjxR8pqxEgqDB5ucJKPY1HvKhi0o6N7QzmLZw/Yiq2vsR0EXuIUk0XIcex+27BUTS/O
KG/uEHaxxHck7n/v7R9ozm9KhlfyF+ibhnLICW7ItdCwPamBAI9ehDaLLyaE9KeL+DLspohzvMNm
H0JN3mJT7kGASzniUtCKTKzzesE7GADLnml94xzk9Y+dSolaiXJjIAsAc2MLrT9oCs+S7mzJZZod
/pEr60apDf6do5P6U9lB7aNcnSlQMW+QkxTEJ52GDZUMO+Hx1vtGJnlhRIhlmNSFDc8N4q+FrfbJ
UUbVb1v4Toc9TKQFxssBC6rafnqBp8RRjye1HnMUdoC6T6YF1Iijn6I4trwJ1lTSta67CKi6Ixl/
G/3IKrnmrUOSTJu/8w93gSpM3fWsOAkXFgk3XR61bLJZYhjxKCzo/xsLmAARkLluNwUUe0/pDOyS
t90a8ySg0o7ZzbobbaA6PRqzHaXLI+SPz+/yoG0WoZPUBUaKG3EDrpYZFMpR5sX4CXJP8jYsbvDo
kzR+dyNsWE8LovRRJa559cAHiD+77OaPzfO8VcSba6a4vKsjO2EoL18sqRkQCBWiDBfYKXIRudAX
K5dko6ZPw8J1VDISCYX2ks4dJs4Tnh2v5B7UNix4tM0taYSzlnpmom7DzQGSqt6cF8h+AW5XPd1N
stz4K0JyK1yRGoXAhAlQRtDMosF0vxcUKr4CIH6I/b5GJN1kKni/tWJeq3sVdsaw8rQnyczYVV2d
IhAeoyYyJu5Klgv8w7h9PYRUkAN1HPyNAYP9qc2PITIGvrXPX1sBxecb1qd+WSUUX7FalF0sSLSD
21QUpPjCKdwfKEiELD6L0Z6M61wdcNyHd3Bry7eM7SSxCc/S98Xf2FoI8AYjg18rmQsXl41vKEjW
qDYuXh4wQdXALl5Q5oxpeNRvKKgBBBjoKxx53YVk3/oFbjq9nHZJS2CF14Izh+aOZtPoh/M5Wcr4
qZ4MM7zYkQHO3QEa1lnssn36nDQ/hIzCY6ExapwXsao6tpnd1FRql/IQK15JbpRbSjB38bXwG3NV
VywkP6P36uFO6oQCgA1bHwudiIS/ANBGMT4Imu+aTWHSNEIwo/ypBZ5IuPspGxGAQ/qDsYpIOiiJ
r20Jhc67l7HY5Z0j/f/fZULUz5qblSR6tyPjHp0orR6Z9jC+C/oeOelf5JV2OuDW3MPwqb+SMSgG
3xnrnbHC3ka3tEwbFnH9tIOJdbKN6cjN95L062q/mh8qmuX4BVd/p5USMKCXV/VacE7nfoHSWD3C
EXXazIUXpRRxMd9tALePdwUU0L2n/WzsXsrVUttRWWc4U2Qi1ItahEwWTHO4jo+7cYNvIIeEmZy8
/WASWG/FaOkkdhHMgJIeTUQwmolVHf6vA1ZBir+9NJ6gjho9j/1zCkncvpsx2DEApI4J484WLBae
q1AtuwR3byBnm5aJD4N0Vr9I21znvyKldFthMRXhZPg+4FA2CBQXoMgeGMW05bUwrkd2gJi1tAWC
7/jCXCumGx29d8BKQV6DYuQq/8jopbq38x4QeWKAFRuSHJ2MROYyXyBOJRZK4eGLPZceLz6TFKmN
CiY4Kru+ggmuY3DrQOYdX+21kZ2gPZO28IjAL9ktx4QH2k+2JCDhhBw2rSI1A3LUQssmvBarR/wU
TK48EIAA+1RwKhWF3C2InFryi4ErV9yRM/1BNYh2yngFbp/CHgGQRblcmD0NUHPvG2ZOeKK6DwiW
5jVwHAZwnrwlA6g6Randw2wcRahPhGmZYR1DU5+dXxMbBp3Zqzo889wAmVXcQg/TtZYu8TyeRe95
M8EcybcRmhTIhuiLPBMneVn50ineA8UArGN5H7DLXer8mJW2K8nW2kDt6JiKcjddF8lcqbQxoxe5
M2OyEsW9vArjpgmHO/Kvqb9NnD1T+iUPUwIGENwSR8ZM5vg2fJAOgTS6huaAK3HqrlJ3vkrv85s7
umwyqGaocAyugcs3AgXccbTwTYQoPE09FxvizcYoPkIKb8qiw43qpjd0qobkWZm5iZWmTO61uZax
USbkzhi8wF9z4zX4J7m4fo2pxvW9/YiIVU7Ff0/FqsiIaxpBh5533bnFDEWj+GlLJBM8UUOt/osG
VHp8uewTlKGyjqPqsHDPXtcXkq/92TROulB6DPrSvBI2o2hSQDyf43OnAHtNCyq7zOSaFdBQHWW5
JAUeGBMoUcIqdJRIVHgEfIQAxGbEUF/op5qcVu2oOl33Qh2UL35fd0JGWebYs/EqA1lwfnJPr4IV
2teYq8f0kJSE57ZdSUOsdbaS23rphZVa6Wi9pqwBxtwZMbx8B9/TdNaq2Dqp8nQpE9nH4uQKpiUF
rM2yGWbFQ1lns9VvQip2eagmZ5DzLIapvHYiSUEZGFszYvdfJzWg7+J8kRKXF4ieC9nA/KCSdLJf
0eHHJ1o3PejNAmlRukm/w4UfdoR5rBbsc/YzkjLwPtg0pkOyAShw0oY2aO18JXISvN/Zm5rhnCJ7
GDV6fdWo211JOgyByEolxRHUxMSLnYMlPkNIcqeCmatYLOVoejJfsVTgP/FemwOvuhPJV8R4v3iA
3Xb23NguwVp63wb8LhFTW0smP1M/jlN6rtQCqQEX5+B6im1/lOLOFtN3IrOnR8QmdaGPpKjo2wS/
QhhEfi/AP0WBfB39OSQ88qn2wHwxt0XSWKLAaciwNh9aVnOkMqvdUBUlUW+YefLwn7/uKKftZ1C3
RryO7QDpzaBZWKMfrWexuEmFrRh5zHCptXmjqe3P1NNsDXlgl90zIW4YKqmcsrPj6RhcgQzSYbvU
MnRqnyTmG54J60Eda8KxQDl3dunf/UY/HZFXlX1oBayCdGKIvg/TGb6E88Oc5k+TrgPm7tOggrN0
5CnNLuqaT5JDtJaI2Z4zKuWswEDKgu0OfiYZcSN40+V6UrtqsNnnQdjH3iGkLyP0sriXnH1uk91T
PJvtPVU9hRX3lQ4+k1E2caykMrmqbpyMv2wUQMsAGLG8tHsoqv4ybzxPR1kXKrZeGaGS5TT52RkL
e7Y/LMA/zDxNNcIyj2SuxQH5kAiDST6CD8Lnfc/Bpa8HaxMS1ZkOa8FFSWjNzlq0mY6OxrfqGdtW
xcm+dh78HzwsfKp/NXyV4KuXm+v0GO3bUmpnVo93DqB71FZc3bAfjmH+Qul198wS9pJ1kWmZXnGW
u8j2XhgMqJgjjswJ1ZV7ztMARPxLXZ2xjGOtZ/OvxGgCzO4Tw5l2PD6fTefuv9nDLnk9TUcvFqG7
bDxS4IYjeELWVvl+mGJfXo2BRoSX/80MCNhCLWi3nDEIsdX0eeJ20IpTMHkR3i5Wc2ctMfB1wVsR
e9IejnGqaUaOnPFGAuvAohJnewDm5mAzWbpZeirrHbIUy0w7hkNNrtc+q0Ve+7MuZeO3ER3mvkCR
BmuLwwyHwjVbGVnv3tXRzvzPFzswe2CqGzqMVTBF26tEeixS3PlRO6SukHuKAVfXGDc0bqW+/SVG
OlQx2NuPpWvEzoqkuG561h831Ez+vERCtKNpn8UxSO0v/kri67GEdam/uYg1EZAp6mteRh9jXkya
Gz9fgaSrlT5hiP24RBkBCK4rJWoKpmeQd7smXxZTDP6gmVAdB219hBC60hJi51yGES/UaW1exl/r
AlcmWb2WgzSmKpyJnQwm96vvqIE6bQZ5xSeCKPPlzTdhRoLdTk5O9tM9Z374wlQ9UPW8+U8ayy+5
C6MGWyHx5hbS9F9c18rp/YdGqlPvsheFnOphbCK5UEINWeqKX72JSpiRtAxh97nTRUvBVAD+fX/X
6Oag+FQOxeOvwUndpL1/g6D+UwhfaAAvMRTGk9Nc4Fqc73C6Tw32DnnSDQE9X3mPfE4OvTKLu2QP
RAkwUli02nMMk5clom/ZNArzspRoeLVhxPmYB4Zc1M73idJtP4t+9nWg5cd7Ie4i1RMHtihYd8vE
pp2pqJuLNhCv+pNXkbVt8TtmEZOLOEysUhImyrgzh3NqB6+9Un12fTi48pA5gTnif4CxDvUmuIhk
Cp1oPlGeaaFH5JMnJjCzYJkbvSWDLdZILZ0hLANYgdA3DoMCv8apjfqqd0E7JgEyCK+a1tLz+IAQ
Aix9qTerWM0o1W4TXYn+Y+aM1EN56jQ5Yryzw6j23I/2hABfBx69D46TTvBD8q8VGJATxnDyPo73
ULKD3w4ZC2335kSJJhs31zwRsHf6GFDt5j6yLdvd1mI18G8lz3MYnGwHc8m2etj2lpsIVPIMYE3L
BDfaox1SxmyUeUNfbrXo0qOdKUBqu1bOgt/TrdD2YO79uXHH7W4lRo5P8kwsJf3kzJi3ZmVhifXI
edBKNLZeko1omTrIgK8zTYl+i/q/FG5eVl6mAMBf/7MoAEugdKwnkRWIE5/G300tHZo5QFgxyrME
+6LxN/NGLAogZ7TDDlCVz/0kNmnfQysjDDtxSaQSpxfDcVR+6l1Zy2ewJoiGPZ49wABPwRQzbQ48
FQDywbB52F+FBRfzS2H57yrGEGx4AlX4FTiG3sA16DmNhfcSzZdN0KNMeCw1MWkv0yzap/KQr/t/
Abp22ZiyPP2giWVv7QvHMtuIJGdnlSZslseWnwBengrLQXdWstyjKQJNDgFOb6lmp/GKG/Kj4v27
WDoBZHKYLLA++pXk9PkNxNUsnEq8ltLtTIqJUBoPVA6NhYhMPCCLGoG2K6xzD1EzURR+ar+LmKb0
fCZewXQQLhZxs9DQtnnbGywICt9JDNpsl/43jqY9HKBmvmhpQXhM1i3LQ18gF2WfzwF1qdcCcyUr
v1JuIO1GxoEg0n1fKC1DOZCNQgbziDxBqfckCAEtMrldjXpPo8Eih+Nxk4AIonmbR2CzN049lyiC
Wl+QC5yVdu/XvSUw3o1j6itcl7y8okxkBNYxA68wRlAbAsLnoZwzYBEUEMtfemGaVHepwMz3tA2g
AwBMASl0szsO2RKavFVc9RjWdGVj64CnoJMRStwVlPubOSSgAgH7rco4HHvSmcXEW+4Ad27/aO8h
pQVZA1Iotu4RexwpAg0Vx86Mv1Qq4s349ssGiZhL4HIWgF91d1tqIDf1X+eRVNII4J8XKjmSehub
F9bq6T2uUYPU2Ieg/9NyqGTM93PJxaxCAldqqrhd/a4jiCZAnXe/NyYJR14bqLf3anTV9gPJ+vHu
GlMES4qdPj1opdJTJd2n0YmfKB6bryVTj4XILoshkyUzSQzmfFaTO7yoIUe/1LD11kZ80GK0fJWH
JPruPwlUOFwSKngzDM7yf4/e/o/zqm+RdZF/PTPL+4waaBHAI+e8hyhpeeFSFJ/7DOBsWYv3gp0B
7EEKR7Gmfvfr4Ue8kCdp4j18s6pnO+9E9vcYbMOZsbPwkqSAxYhoj+dNAivJqeSO/7jcSUFbszZn
cwXr/Ff9XS7SqX/ml+xjpxuysxZ/Qg/At9+uttvESPhAWPxeyTYxd9rcmvSkyTRWfg66zd3QNhaE
EbNrIj7XZegudpK9c/yAf1J4NxLVn+5W36+whW+9PsJG2qG/8eiiI4N726Lwu1UxUzOJEFt4SzjF
gmzbDPmZrPyOKJUgsrh9uLrc0/D2QzDdE5D+SOTLkdIoj9j+3KCgTwXeCPRkbdaYkExhOSl9S1Fc
ESBDm4ouriZu2R1mjRdVpkcNaXhWlyUw/ZdcHyIUdDvF2DWrn9usxrHkZHWD14Vwg4EGnmtqtnRJ
NnxvqKSl2KwVl2Hpa8zn1uEI1pW+5FTXl1aAYQqxeQNmwEPHzmP6VDzLwOHjnuu0bvAY697oRp1m
wYpojfaBd6J6R4AnrbvvIh+Y3FMZJmHiFWSc8A7Nhvn8cBi/eULYN3uT0dRh+ZQTtaj6OyWVgUW9
JvN6OgLGVMBeV2gnzmzPZhlZk3oyh8eEuz3OPaK9vIAsTdfTwG0x/uDBN3E9XqYKCEXDSTlAE3V1
yXdmmlAcUn7uI5wMtEU40w60myBM/cymf6fiH/7q6Yzn04f+13f8FmvNv9F1sODan+t4/9euOd/G
okRFbxzXqvgwOeHWt6o5X2aexRBU5ZpGzgxB9XEV/3SqIqy6eBTXET8HxRLfrVd/A01gmN5OI1AL
rRYADGUrsJc67Q3UxaSBBlwdTPikNdX3VNcfjD6m2SlJmZdtu4LKpBpqOtWf1Imq6ym/QugLzxee
1BFpi/RMDM2ZSNTEdKOnbbWRgRxW90hwpb65zYOEwGTN/miQlSTIKiW7nBNALYKz/wgCJxaGk0UV
AN4sTGFkXRgsSx5VKnH1RyiSl9k8bK7Io9jxMW4L8nGEwBRtW3cMurMyXfSl/QqjXEeASyyKB014
crsF64EesCwweGhblXRld7DmcQtue/+0NoUxQBB8EEHQCsnqSuL0wENIxvDuHOPipiOetqyHACz9
uLGAnvOOZzsEqbX6jZk4/Vt2TuE85QOM3JyIendgM/D0qUWV2BfqnG4okNNDfgFGP6o239riKnrv
B9J8wtL9C9vLUDWzYO+d/YGpQ5CHmTbUqKbomO9oWd4TEX2N8t4SCXZjbek5rxZnARYEpQzT+vvw
ZquYS2Ym5OHoGGY/ADCds9+CGbff5BrwNxnSAMGkXaErgErmT9AHeubdQXhMnXwsIAiQgYFNWETI
FbAaWJe/HIHlf5/90icyMf/R9TUBhxee/rOo5noujWPt1VW6nIqVzsROQemnZxwvVX9+Ht0CW6q0
QnGaz33Ukp70k/cPbFBtZ2CSHXKGCZygeCwbM7jSZ8OQE2gYdQGVhXTNrNLpLD0ioKqC0vvD/6x/
wlEdPuF3Sn9/FCvhqp++PBhsdFMOfdbxRrgMKw1xjzSQoTYJz1idnRGHYikxFfQ/SU+ALGNQUUo+
dmHk7nHWV0MT9hgOXgelSEo4+tk78wK6OITLdyIxYI962M3dcsyfUyLZbolRhdoQZKe+AQ4Ek91h
jgvXN0LYSTIJ8jSpmGXgqpVksgke9mtRoaFccDdXXyAtGFhts8zc3hgMB3FPwbe9yno0+GD1yem9
6jB3/ioHpNli5cE+eVfjwpAD8V7q1qnNpa5HDwwyp/WBeaMTHFqQOoGSqogFaFg/Oq+zJTfKlLtn
jeRQom5B7LaaGppmI7Kl3GIsTLYUWniQEYilqRA4Jmmlajr1aCcmr3IQLm8qeca36MMPv4POX0QV
8Hp26QwldwGYTweI5/RjpQxEAlFrGScYdd2QTZMJa783rer9bI69RLE88gX7qI6D2423Un+/ZlB8
YfGXuGT+Id1KXKl2xDgJBowEfpxSNEBC1Js1PHJ+74Kx1XPfaBhZG/VBjziZUwYUmeexEuLAwzQs
WEnEb5rdZaAogXu+jKFOzXnoudnsxqbMw+xAizjzLUtfkzgTexj5/wApub6HhdO76dgibfVHJxUJ
HunthIt4ZWTJGnLXEYuAXjEabRtl1a6zyLeFDubQPtYH7WU3Koka/7vjA153QzcTby/mqYXm1jej
79VChBs5loVJDyiJES0Zd1f+fGzmuu0CE80m6gzVwblOdKCZOW4caEIaPYKX+L1R6loxBi7zs3wT
OcVOAQWsigv3BLBUJ6PvsVgdXaJDex7KccuO1EtutVYw3SYvKXZX776fmaFxpOYjjUYfKwkCIC21
Pf+yklo6r/ETzRSY7NMEh4cwkznfTxvoynZHsvdcgdFkEBacdqWT3/G96nQ4Z7c7akzhaf1nGJL/
Ct9zgo/Z4umBUVJcSoms7K7lNT7RFbQ+HVwhXMyBwrBMSquIUnRV3KwnsWHtNeaIR13ksrpKSDhf
7IAgChYY8ndVx0xnnnl5tkE1H0byBPsZbBlOM+mhfGDYWYDPLjXARSMXrY6uWeaFmTDK7WbGSTGT
z3b6MPk0Cjh+JfYcpUfaOWlSkWtmAkR8MvWayhlU7Ea3UhsET0t6r4BEkIJI+GcrydvI0Qz66ViJ
24AvTj6TjO3j8v/5+Sof8XK/Ow3lHfS9+iD+I8kTI3uaK/Z+g19aNuVkiT2xFA2BoPScHfI6L0h2
c1ITNnOgXS43DZ3mKlbd+72h/CazKUG18+IUKBusKUvZF47pjaU6oqu24iUmwmHxeUrcUycwQUKZ
DfpKO18+vr7YF79Y1iD//IWVaPbnl6baQxW7PEU/x0SohtxECB7sDi/Bo8QJX8B5fN5NLnxkkoxy
1j8/W9a3t7O1T89jE031T1qc4U5n+5W0mKokn8QIOi8uGpdrDaKlYP0l/Kj1E0h9v44TEKHTq5p4
gaNu7VWY4OkDKesDn5pamHiI+8g+O6KvprH6hMLDPVrTHUhKPvF/irmAi3Ec/XgGSOAYYBNcMcLg
kS/HuGc4SS0Fkc811Nn3AnF4w+CZvm4FKsOlC29F7LSDPa/2Mf0yj3FZJQZ9iUiOW/X1MgrwpAkP
rL4w1i26oXtNs/GqSqjNY9jXpNonca34/92sxLeuUJbnQ/D6eSt0F0e5AQ+LH3mH+wr/RnS2UULF
AhIibYjtdhfvl/48LG2W7Ep1rbxHvANTTQzPHs/V4kzvOdGEU3YA6G1hxgm/ujnn4ezqC0O4Pdi1
jVPtR3qQ4gvaCOctwtvT2XRHQFlJvLg9Eq8X8AgKJtYmHAeUzZCMBRY8EDx1uBb1X3HPWVbycc9s
3aRhpMeLR8tMPewWdafBnBjrbL/hdCFpoWR9W2qu+4oRZZ8xYtJGWXSP5zTN/nzoQxfWU0eKAhx4
3ikiJwASVMlo/icufOFAgcChZqOyHu3n1alXGciDrfwteZ4DdhlR1QRPbB+TFU6ifC2+iy9d9XlL
NMVbNpo7YKjZNV8G7qvwHzXo8syDbgCbkj/YIFcDKXFmalKKXGaFQyUc+tOBaWJ3wrMkxJNtMv13
JAOzg+veNZ4kzqO7NCQVlpZR80p4aHFWvgyOrXf+jdL1/YKuPOY/6hyLp81xdL9rsIrHtDRZeurC
vUdpAsEkc5cuqXkL8HPCw6WkSahfze+Fbts7YjbX3rUmxRw/+6Ob843t9hLFGH13q4YBQPOrNwqJ
wSEg6BTgUuY8C7XpMw+t92qaCs3lb3RH87rbFFh+7CtfAJwJ04Bmzeam1TiLq7bLkJ/53t0R/s5z
NSN2+aTyllGM20p4lgaCtyMHuzw0VDpp+A95qEi6umHvv7jS2aL2QMcTCGLaut3qSFzrXn/Q4kK5
YaRDqscL3tTTYY6Yn+jhcDOTEkMErg+4GmREnCYyM6CYxLPOyEDxwRs8h04TLDEkZPv7oQ99YDz2
q/RAAGOCwGoouN3m0bo8k0hOEKuXPyU06kGDRNaQAovtd9oPF+PcCEZvkHe1Q468fQF+5bNbdqY+
J23YpeISpDPE/xCrr/lD5foY7mUIh3PuMmN9nT0Vaup/i72MPZCJOSGCcaRvdgyIvB4PP1+o0v0m
CDLf1Sd4SUQN1dxhf3edr+TC0SidPtvA3RXg696Oxwm/6SrjfgPePiSN85PzvpJA30Pax8k/E896
VdBC4vyYxdwe1sda1L1rErkEKowQlrmDGQsykuSa+nR/ZJ/eYytgRKi8VlClhYj48/BQEegyZ1xK
UJ7VLeEeONqHAWg2+JL5BXuImtPm+8U/8PT1CFsp36tWjRnM7y78ryh+bwUDW06ZJUKmcnQ20BjT
kUotrRuOGNW3jYjvVLhjfxw4hT+mQX+kP8Z9RJswS4K4FIIiGvXaxiQLTWzqmUr1bNEA/vMvWAl2
MvqIl4sAQO6bkz6+OScEyQ6wm42GLoSGQ3DnDIgPmFYLeE2XDXPWcNR0mrwwXlvyfCqudLoOhuNU
2zXc4J5JBHzSpCpatq7QsUjVDNdJN2mdhYhuadvpR5gghl65EZEw04QaRHM2kCcbNY49rfX9gBhb
wukJrtJXn5VjB+LwpkOy8p5wwZs9IkVyUSfhpy8To1rHDXI5HgHAysBWOvLoFb8YjLuioQvcnrUI
S+ZVu0SirNyp3XIATmj+Q4cx3eWd7gifS35aDdegCo8Oysr6Nm6lg8J7mRptnJPuUXknqeaWe+97
woxkd2Q595qQR/DOt3Tyuau0wIs1fYFO0W2IEaU9iOZFT3xWTqwUpPCMVrvw1U3IIgvh4s0STCjj
A9UMj8/rv+csF0KQpz/yMXV4aYB8MYm47cvQTDIH2tS+Hz2T6aYtzGK2zUGoTg4ELSFz+WJWTnbX
VKp4luEkNoqPmEoaZKpdrfNZwcG30RmnbJc7f7pPHzLgZIBRubUJrIbiPrO8jxiTeoZ1o0gnjIJI
un4UJU42E7HJ7ds06hye3qNi5cIWBf95kZCgq/0u3kpHpZ6XE67vnhxAXb4D8tGbOZcBuM3AXbBw
BbrwHDBFGkrCoeINd8dimofRKU78PPd9aBYW+oOQdC5A86+pL0GXAIkNf7OTucdNTUHhkgR9zc/E
/sHHfKLoZ6vebEDSIwA7cucgBxFXMKjcWzjUr7rhrX8wD0TPE+EJftNucxP0C+CUbVBoyK3ZNDBa
oBLsigFsjzInmohyObmZ40hQaK7Bje0o6gNb6fTl8DHw1LCJGomL5/ISvXQhRP3CGZDt1JY9e+S2
0drHYJqIcQ3S2lok5V9rDKwxuHuGMf0qYDnaG2VV9ZkORzOBhFSlGcKpuW8V3+Wi7Wg54RMCfKTr
7wbSlAdB9J4BxUuVNVJGEWWC6Q55fG0TBjDryOenjUyrUR4WrZsJ7VPPESpsKCLpH5Y9zSnzXpEV
lIf+ySPDt4bDtgc7b4/a7h0u9oKc7Os06JQN9GxOBgVAzeq1PCWYLOwSC4068ztzm+XNNWXnaoli
/+/moPR5TZyjvDzOOOb2KziRVINhTRoYRhNstXI1PKoC34kxOTvo85x3CmMCkCEyjQgjQhdjvduj
A6oRnSVpDnDiiH+s+ROnufVuhdh/Jpdxm/oSMvKe/uyNNoJ+SP+rN1EhgB30w6IZqvq4CDIMP6gU
WCb1T2MLpeeI9AL1rN736kq78H9ufv86AQOIqJ8MN4RGKvsVWJiaTGJlvZ3EQjGc/oDoXN5ROG3H
LOKjsRfWpf2aCaFYiXE9haGXFRkiJJdxn+AODWmsbdvhtOEVIqMNlTqVecqQRTKnt4GOEGId2h1/
Q+Jl9kJeKJ9rEs5Ovq0bhncYKZG8unXpjsUbmVs7WKGLsd/DQJ1kBg45+dxmp0KL0YjVH/P2vmRC
3Xt5+fcChTJ28rzfFjlYh9HO0mk12Abq938y3tGdRa/PHxpVVEqnQCPOQ44H+M3DS0YaX4gyKzjn
zGYvgxkph4l6cn3taxY21gfh2ljd6QpB+Om4Z4cpMFdbft1p+a9wLJUp74l2xE1re1HVtvMdNspx
TasJr0u7mpUka8mK2z4ihwRPl/nob4RjcnGsSrdI59+OYfBhWZVprst+5V8jslQBoQKsb24KGBFT
MGnAo889J4yuOPXKCVx/89Dsx5lV7SBH2zQJqVcWu84fhKd/iVyxI29BBrd+DEeiP6+sLoVGW4G+
KOVi+IRgoUOnap7njqVXjTDjoalybflGFE4CZjLsR4T0J1rYcskaO5tzZe1VgZkYR8Qv4FPddaeQ
fw0vGF/Kfw2FuiubbPsnnmfKj3xG9tRv+aONU230TDL7q92MGiqVvu5GpoMUU8OfsrFYLS/ZAnqU
yBPi/Kp0J+N00q0TfYRGbW7jkT23Eb5ITgSiDz6H3sp29QwwcfpVn1VvusRyFPJazHgtN8vYurk+
dqIaDP2Fs5iSP6Orl67FO7LTBPQtvYYlF0BqoDWffGb4lTFqt0ziMgbOwnwoy+NbGaVdRewq18CC
tiu4QfCty+i+TJ0UTotZxqT8W+yWBE2VwzGgp8F5x+IKXDsFCgzMWXu3RwBGpgz9nfyp1lI0yeN6
Tx9G4wyvTaLLPirLMct88AsmVh4voBfTbrAEDDDU1VRJoisP674Kt2YmEwZyoYeNRxEGG6q0mXRy
12bicsKjNUg1xXhzDyELI9yC6UqLUX5CggATOy8IRLz087/NFzdfWSwzQ0+KIhHsw/Fc7Q5AZDjY
8njoPM9Tm0WrwYMcbuFnl68MJuhQiwLsLV1O4b7TsvPM3nAFPDGvTeU/yCQIYkL+tSUrynfCbaLz
EXb/48JR69r9EaldjzsIqtHRSrFlGBcFY5n/DQiheN9mZ7AW1U6uYOMWqtt9rE5DHNV3g5OnXD5u
zoQZtjzOAalMNy6GxGKVZSk0rZKhafBYBemRg/YH099zYETUk2AWS8SRuc88g2To60lIL8maUbiK
M2kevOqx4alK2XCEJ1hSuzYy97Y/4/yvUMBl7JNRHuvETX/Vqw83iyo0K9YLosSetZtCC+lBc1I3
amCJHrx2Z1vizl5O8jEWLWYTXdcWaw4LLoZjiNPyYr2SPl1CiUfYanAzKJu7EAuvb1c1TwRu8XD6
DbWA1AsE3TaTy/RarpHTlfBQlKX+IyIev/V83nfy9G8myendWK7zAkpK9RMBF6hIKf1mKCZKovZH
V+DoIcXXD33CjQbBcUumyOiPWpcLOx8gix/EQmmwriAb8ddR5HnTlEq04W6GOAYrPeRR4gqcfUIg
H9kctULx407UJsBh/WDhJD5VyrTOx5dmzSh+vIcKSumnEqy1hy1wHbIZFiHRAtBdXXYeNbsB90x7
KjldIVx9IkWE9q7uPOm1EJ9D3DJX1fndCs9Cn6+f6QV1RUuzm7MJfd+27s+zYRP5t3wEDNCRZ+oH
oWy1NVUaudGiB+6BUrBhmluDHeHyM+E9EX9Et38uj9mlfa+crlTjP2IFfc92EFuj+Fw49m5OC4r4
55LOt8CAa8l/EwfMGzE7rAKmP3nVWq/bHfHs9PpjPukdJYBGKkcw2nFliPJ7gIPNaBKiFpsxx6hZ
xJxbuxnSyRmuTuxaVyx7sG2eNk6rHCvbkVYKiWxOOFpb0duUItlKWimuR/q/QFymg0SpkhwC2wJN
JsGEHfXhAOd5cPW5fPQaDC0vSonjbSbK58hoH8dAv4nVPWSfYIxI+j2Dos13b9EqksBeEfYSn4+k
rNvoq6aQH7q9c+sA4A+vvKF24eSK/eqJDYyc2iwhDm2zXONFj40OyXLExrqt3V0hZpRItwJHWC5i
lQUOq4Dx+AD2qNmypnngFZrIyRYdofVYwJuvTbYxfmfXTTWYsqfuMfSiTwJfBEiWs90PGFCCzT+H
CoTC6EJkBev2miGFOk6NQM4C97wCKP+qPiATK90kYS5qkRgTmXgTzcWbNt8B6D1SuSTDbtkyT7rE
cLbzgM2nq3qelCGm/sHRJiF1vUS/+sRAsnlmcefaCu3yWMnrh5k1F6gJelSZmNNZk55bFhQ+dKyW
BCLqjepoLZyAX0SlQsYjimrqLzWJbiCuMD62Va8g9NECneIfPA1enksePp3/KxpnjEEflLzVnnOJ
I2kfKoF3h2nY1PIP61Q0/Gp6puU4LMKP2y7ksBTRKAVcxqsJzUM5qBh+AI3wUTZul8Q6KY0UlVCJ
h7VjEV4JFYttDF0wX7UVWm88BMWt0yleZdUdK0ZstqDFcwxkLDI9qlQNcTMThOdcriCK1u5jzOz7
Z2VVjeIBKpeE4PL9mel1ZskcLexjBE8/kqeqys0CBeu72caTmycahr6deETtJCUqrh8Chgtq2+bG
xJa0jeoGZjwO0dzPIcstNcLtYkkfEYgXuGm0silH5O91tPdNTyghmYnc46FMAHg8AVtYy6MKUEhe
lomi1A9EO2Ga7DIeUpywg08uA//s2inQMJFC8VC/xZiyOVTYFRo0rpL/FJbK8+JZJ5H3j2Qg/KcD
j+0YLGuYIhVdsTyrtwBcWZ5yH1h+61zV//uhGtQVUqwVd3JiMGkUsw+U4JDkXh+L85hb0fowIMQw
TgvJFpBcWGkiV9WrYwl6h53p2mN8kQgh1Wo1J6V4Q6m2L/qNtYt0BOdhRCjcnPnAYwrIwHvhQRs7
U2nFT+HGxXBDFkunWbMQyGYwNf/yZM7biWrTUSeCIVQKG0YTSOZbS/5PNFuZz6pdaW4UQ4jC4QG7
fhsDitwEwO1ievOV+mHOg4079M4rpMkG+elvtCWHtGz5xwRLYnKlfbc39Uphlk3IyVgR+z/KUH82
kXfdUgsIw0RNG5kLvGrrQ1XWR1RqSoeZn/85IAgglxCPOPlzKOBurdYZ68osqHMZ3FZA03e7qegD
JPgMaP5jQ+EQgDr2DrVFwpqEZgJ+udUYEYloUPSNUVtjw621UJhm82uphdoRyXequNPMHsE6wuco
8odIBBeSiX6771Lsqf+zn5CEt9tJr71+IzLsN6x8muxFEYVfIeSqt/WtdQQ/Du7BoQwIxBqH2UA3
tpKcKMcMqKCx386e8aBQxz1Oyg3dsmWSYinOxYY6y3MeRFTNxXQFFp+OUy9onUDXap5VTXMHrOkB
tGo/N8eRF58A6uViGmnhsZ88vnOD1zbQIhbOfnW+IHzyNK7ViIdQ9RvxTiELHhZm+nSVK68THgms
ZN5kYsFvi19FdXyfMRq3+Rb165NscASOMMDeVm998QXCVpKVyUubuUsPlTyXJteCa2nu6fiefeK7
I95Dg7Q+VO0dV6d7XQiB+YJQ7Rjp7+yiB3JfwRws5l6mlx0ajDAKYXghrsZ8atl6ibM0G2D1PBZ1
CnlTcOeM/jPoPRuhiJGXPha1fnZsWoOFWRYbCJu4pvSyAlRN537/M2bjIhH9tgFQ/S22fXAypISM
r12s/Q17UYfkeMeH4nDx3AqkO7JURa+D7QQHMH+DjqZRyiTJAL0NPdMtb4gLgP636yg77HP2hVXO
HCUuqFjSJ+e7F/ChF/q77fhHAUTEa06pehxGUfTcRYOXvo6BbWeCE7r/IIIl1zsNtppbSkQrOaCB
THVkdfUsMQ+U9bkEFDKchhdTn6iYJ/QmoRej+lWJqF50Q5vZEiSFT6GxSUNoNRphcDa4GZ1I3zK+
ATNnBSO4PksO07VwkA/NEKvx9hL/sN5PlaqfUoaTmJbWOYYQiS+VDMJVUtJOXSP1nTlCiBTLcw8i
VKG5h2OZwpf4tBX0p1b88t0AQKDPjrkm9Jtc6iBbGDZM8dmVIBHf/sUMXZL5HZdXfsJIoLck4MrR
VHKUB/uqIdtHvpI0+oZHA1ruoO5rH1YH2jFMGzzKOzNYaOer75BdqJCBobvOxqjsvhZYZ0yVT6M/
YTqbTXQo58Uh4J7hfGOVjXabms9HgbjPSgADxTyi5v/RWMGrqmdI/j2jw8dvtFKjVhp2Ix/mZbDT
7Glx5fvQ+q2APJUNqsAzuqxEaytpRQvfYZxWE15PM8edHyOToxwJA/RbZJQgOekkJNBfuEfK8ASC
8cQtlmqqJzRKfRvAMW9IP+bZyl1OtgOyOed5D9YmF7kuqDe7MKRgzxcZsVghBKZwyTsZNrNzcn7b
/sqDHWrkgZzGv1FNDRqXSuhvvSvi23btbG6U3fx0Gmh35rgxhzq6kZxNyszG9dWeFiFw29YybipF
kBdyjWdDK5QbLzf4u/JEny29niVMTirhdHIdBPsIKb+eABN8QDBjMXpsBJtr4iceKhpdlcIa4yPy
12581h5mbiQxXqfQ6hHdpChJgVPy6/KA6wwKSqh9GqgXCwt6D9UVDMOzKq86FMwgOfEWJ/BjjmNk
g87aL1CBWExGObzZ15+AHCG1MEWT4Oaa3hLj2TUrvLae2z7fVChEj5aKpyEHFYPl3s+oCSPwZpAL
8h4RyhaiUIF5HX1jV652uJnYCxRsxOrxWBYmC3JuS32Wwz4DJ+PGv+bqpHFnDCCe6YCrbp5L/jxR
vgq+G+8yMbzF8jqLhulKdm8DBadLkqSpwE35pfyfBSqLDte4EDG7DqOxXmQOH+lLGXRz3KKdMG66
qN6mx8ubP/OjUzkxlCt0L1umNm6+cnl7MoIKOM1BX4SecTh8UqPCOPyBpJa2aZ+Z164nM9ApO80N
gkpc/7/I6PWe1xgdQRM7zwJ9HwxyLKQZF9NAP+RQas++OiffMiRvxgSkXXYmMvEMlEmiv7n7oiON
9sRqXaQl+YSUabmvbPfAFAdlXt8Q+rW+08EgAUiKBJ7SuWmFGjoSHw2vZFSxi8XYcAIOTva/kxix
712L6XVQu309yz+Uk5fItzqUXbg/xDVF66AwawQOkku0DhJCShIxJunZU5DOqp4iqHtgISBFYzuU
fXtWD5zhkVU4AKTaWHe9DjgSPgks/5KSYmSZo9HgrKvVrzcCgzYyh5rP3FGmHIPrDr/kQ8zp+Q/J
ab7+tDLiD08/ZuqDF1cUw/4tzNRo17frCKkL0Lb++cjFOG4vdsw8ObqxcRk2CefHXzdgCGMp1QH8
eTdKfNg3MBxQty5tFc362iaZTjlGDSa634RzJ0ETvO/VorG48A66ZrYEa+7aGUvd/ptmOppotTL1
jlcq4RS0KPt/R9aTvQCbailFDrI0QVpLTlFte7OzJKwbi+Kj5uu4OjGCePqUgIAnbFnnemEkhLYT
tSV8tS8nh2GJICuExfzU9Lu9OYDZvtDzRBVDCw9WfkBF4fQ4YwohCVqNz6TnvRJWUfv3k3pz3aTu
GddmLcA395BhRpXqiHjL5Xyo5xDtjDoKNY8AnQIgu1P3eTK4BCGazuWjTMRnQ1LDMc8HFq1lOO9t
xEKUPKQHDlmpBJg7Idzb6pGyCgH1N8sPIvWtsJnsG7tS+6nvLr6ezvtoPPtkE+X18yIa0x25AMAy
+ND7oXSyoAvkjpDLVhYa/bpdtSgUvEz8LfUfkWcP/GxKYVqr7pz7KrFR3uWhqqOIEnweMG/FkZRR
m3P8Qv0vuHgw8fu5vY4/Lu+WzffGAa9TscZa0HudM2RPYbKKZ3XbX21ayzCP6wGgsgPz/SHOnMXD
tTf5IhWE2NckFwDxstEchPqgj4o9gi/Cd4oWXRqx42BtowgwbqmWq454xe4kSLGqJqG00seRYkds
QRuKOACB0PvncTZ4g6if334wjfKXzbwaxngqdPyEXf16A9BwBHkoA/m0ee4HP/miydHbxpbqThGK
4r7rB3INza71snGE3PTgRgXll4NhHQrX7YdYtaF1pTWJOjQdO6Jd4/qDGD82LSbse1baKygDfu2P
mwmY/t7xErgG9htoVIEFu1PCfpjZB9/nMHMWQAYBLzU/NvGivpmr/iOe7mX3JUunlbVEVhA9or0M
4o9P3t+DWtwyGcPvtY9nhVTtCxfUbnLfiy6Hd36GLW+5kWLz13ou1kz37Bx0NL3EAhDIxeDVoj6H
X9q16gSOuE+9ZnFQIx44h7HQ2GgN0Q+uzuBU8C4uaQEZZL7tEPXxuQZWqoj3398LqO246B/fXasz
3IjcFbm/D3l/RmUs1MhDCKld2nL/LVqHydvhCkXCLDrNGT2iYUzWSwcj/2wKiczUr7InnIDj+Fon
ZxGfw1RYmSLwGH6ooJuI9aMwFKfunsR+ANDDgH9+gieOZYBp5kYhL27kscVjoLaL3fM2SIHHg58o
PIEmQGH6qW+OJEP7Mgjo3Sx6pp2r3D3Vmzwb3ohzBgzqTqB1JLk19OIYIw8C2QnbVwjucTy9tnd0
eUEDLtJHWqqpENq9EgRHcIm+itV0H161MFKUpQ/7g+m8q62stB0rwQWNk6N+VgJ+G2+NjcFeNZP6
B7XHQ+e5GmHdzmGPu2wA+pqJafxAnmeB4tvtgrSDHLwk2iPpSfq//1M/D7vOK+KXOc3sc6tgzemC
9EHjCmBCHj+fkbRHSo1a4DeNrn6ZfloZ1RNROackO9KuKB9yuw6MUBri4ED0O9Y/ZvyhivHqoDH/
p1eMomrsGlIFjDLjMjH+QIGXsgY35Lq5dm/yymKpOMrKGfrvmWHN9AJoXVITjxoCuu8E1FJ3qTdN
FaAYJ19Na/O48mQrXJvAOOU4CqPTCSBpZ66xlar72Hh/49uMc010znul23UDqYVNHVxl/rUM1ofR
CdqOQEudZrauCGxGFTYvyJWUUVAfsrF4kIbzwNVHML1XerHLMlX7XOG/Iq6bqDmIJl75b/eGMmJ3
Y4/ciUN6enhchUmR4wsILaTcPHjrjky42k5TqUINA/gT5NC/zXnp6iWMVZUp8KRcj3mr0D4TX7as
M/8Wsc8zE2d4KE3vDMaJHEQ8fdWjHXeX3CeV0mE1oy2Ql+4LKRNLz7TCYJoDg9FUe2+soiN8CThv
X+3dIBNVaMkzEwQ4Co3U/LV9Zi864QbtOwvvyCLUQM5WS1WYv9IdGGpoQlXge36nffEo4U9e1Nsu
Tp5C8IFhgI6NKaBmitcBnCR/hHoYwNHT17TipET6q5EXyUk+OJUalGGwktAt/RNFO2BCd15D0CcP
5wke6i8Ailt52oWUhkkRs0ycQxd0ifk41OPDrQhZfeZU8SPCUtfJd6TM3oS5I/uJn9X3qlNApLBc
WDzP1y9IHr2uq8EqkXabnvv225Omd/xN9mD1g+4My/B7s42nMOhK0RnN3sVb8b4Umpmn+voV3Vwf
WrKLKKvgcGz9h09ZBxTVsACekVbyef+aUX6kYFxP9pEGlv+VpPr6Lpk41FlcDhEzD24qHuQ6iNFv
DLloWDoqyqV1+4xp0tuY8HPPc7/uGa/ACcAxJSPd9QiZUdUEK9c1dxNUZBtx48Qg3/vOIBQ0+JFT
uhh4yp3lB1VdbmLM/Fv+iTaPq4taqmoExdCnvJjYaI1Ka06OfovMpVk1Dxg/i3ln1GkcLdP90Ak5
kdKqlpnmUaI02NOrIFEY/wgbPYMX7S0G+BPPbxFRN3xd2O5QheWEwRPPbPF9ZebtKA9k80Ls3PPc
wYFrPmN/7LqGixS5tqf0k4mkVbP/AOoirNWdLDNAsSm8n7/+UGVhxy7+zRRoZTANljGmdkLT+16Q
+G14HxwHpWUAxzLCjhZWH3PYsJuqoeTNA4P8pfl0V61T4p83TgPcGdsb+2rjeZDTj4T1YqUWdGSE
TDCpjoJBk4RwFHh1BTOfHMkwkw+uVkHZjdOEuXyHPaBgmzTg8CCYV1qxfyLFoAf1slp9808/JqyH
ftOlQaik17vVWd6zkcab6LAn6Sdo17Vcobwl4V3vMGb6qLazoao2ZsWGOSke9BQdeuFD+4mBg/k1
/4pcMlCkz/GKFqGKwnWm31zZUzsw7oGUEkB1g+T0BZa1/R9uBfBqPVAw77051XHm6S8LnYmOkr44
qG/lSY3FUirz1vCPHzC2dYMVbvgdipcq7ElB0CWur0RJgZUdUyqNk5yfI4unHXqYlhn843JuMIHk
BBwFQji6d8spLxa5sUPLyanq9boCrD8GZN9yj+0GeeWfEgyUM/rqx52qcCra6+/jEEqZuMaZJOub
a8N5OQsdo5QkEMEKOBbF2X0mAEro2E7eTHzQhAmGbVQzfB6QV02hRRXWJpCN8/NC8L+McKow7Dpg
WPB71AqB8t/jMp2RFZ+aLUplYuWxRjxydwTv66VlVjnu3Snhpk0Xujrfz4dkvoAO9ADFs2hT8yVM
WaRqLwu0PXhrsptBQ/DI7iHSNDKqQb8ag1vfeQStYT11i61B+bKO98NDbpU+Md4Bn8/KzXYXpIxt
eRel32oQIEbYpr0XG0352c6Gr2j9TRoEB1Mnd9A7fsbQEqj10DFH8kFWYxqnRDkVeTG1lpPWCJ5d
Z9NpPQgkQ31jFf1kwE4hkyataeD2xchR9UhrCmq4aOEqixstL2/jEYaHq5iW3uqxobmgsqFatZHr
xwDuPYlzOGGKQFVCdUqMDtJzfaHxim3CwAJFUdk7nIbOhfVbUAq0hl/16uc6m9lZqt1LwbT78W6M
ANvsHsvA9lUHW7CEa+n3YtMHGvpeA/iXdYd3rx4QbRn3Md+IJledErP/2Rw8A/ZbsVLdUUQ4kV8I
NX0CiOB/jgcKyr3FVjuKB/2zETGUii9M6VJQi9Hi2n6uWUGKwYtnLnkPQW8V0BmNDxrRvx3OiULQ
IcAFsnhWbrY/krEHTWYRxx1hJ+HgiUsDQ58JMKcftUuAWe/dO/HYA8jH4r4aLVbSjDj3gT1Qe0K6
oAiFUQ0ORB8xL62GrDGwj7mxf32kqyWXn0Fj5MD4tpLsOSEN2L2poZdtyp7MsK/e0kBqyPQ5YIjh
/mcplUEaVb0g+Zjc/FgVxVGGsZpPGda/i9aYvfbW/uukKKd5n0ds6AOCYNT5pf11x63cfwJgYGOk
NMhRpFnluq0+DW5+EUw2zYcJPxxPPWZR9FEtdKNTyV3Zbaz64DjZNk9ln07VSDp2YWOnC14DcxSp
cBSRsZYAD5KPkXV0gPUJE7TjURw9qAscIbOTH3ReY4ApaFsBDHQoHhANM/5PbUI9gLs/D/VIHJZo
rHt10uH59TAMcoHdEcEqx4LsQcGBiihHSnzJ+7j0LcP9OXBOesICohNCHSKz0Js1qr1FTRfM3P5v
xpKm44qXgOg9icCr09G/OE3C6c+HqgM25dd5n8sb1HpHavEKq7rHJF+2Pm6oIFl+6xgl6h+BHZpS
twNHIVFDKzr3aycKmdNVcVZCte47Af75lDGkZyxt3Kh9WS0ob6iPoRnpGsF6cJlkGaNh/o5+axcD
F0AasYaM9vVic9ofC4h36Em+ymt3c4d/TTQ4Lw08teKq2DfmHir4fXxMiL2Gm80I4x58Ek8SzAeA
ymccylE0XakSa/MfwGElup5rfc1ZaF7dClXYBf9A3n8xfcvqz689ivTuEYHy0D1ugiVyFTvJS77Y
mAlxn84EcyFeusnEk4YM7P44MBdIRkec35/EmXrAB2hH921BTiTHx5CkhCV+IbUP0Y5plpfcm9D3
sYtlGNCJsnH4CQ9KwDgkhqQFA47AyVcB2SOhXkj1FpHlP57oGICBAo3jLUee8JmYM/i7YVtW6ghW
owpgT30+oGLlt1sDDUKmnH18oZiE0Xz6YEPGZADc3W7t/InQXWwAXVVhmw0p/Ne1QkWrKvj01Qqx
MUoIG6STCwmJ3hVSTSPBd3SybwH3BRX1OI1F0p0nQtTRxwPEqUh2BXq/v5bbhlHxbPpUObt5b05B
8WP6dQJtgyyuaqKerX7K6KsSTJdhM5qzUlCqgUA3ul3ftXEXyhdftpobv9z/1j6HIaKy0IxXxFUJ
Z2+EVp5s6tY81+h5ZvlLhUvF6inFkxR9tVShoYfF2DrK7SUh3J2B8hvnI8jDtzln4AzR8LmcOKco
np4rtTfy8AjNAl6tS0hctPUZhyQD6gL1ULmPGtxDMk0Z98WgT0SJ37zk3VjAXQjVlfS7ujxakQGk
IBXy5hR2J0nCYlU629/UylhAYcSwxZno81swlQCxe0NAxpMfuYEnKwkWNJ+KYmkxrErrhgwzQEyj
tzfc63UvIoAZ8s5eTZDY9rOxaflkB0FidnCEHwLs5ylRyhrxsEQNGzGdrj4uIiu1GzbsePyZCdvL
1bi4++II+zbzU79inmjQU0dMJh+6J/38e47Vy+FgKRiclKB96yWswGRUGhhZKQZfm8Gn8O1TW/gF
VG9g6qNJvQc0yVTa0VvRIs0KYmIporayUv5XX82sW2eGuuaOioIk2SQMONhXfRfczgiCghMknBZV
VU3JJoH/yhK08inU7mg7f5MOTN5SvoSJpKA6yFmetc+qGS/QQdVUUAWfWQ2CujQVFvGuxvu8tZd/
Q1FQhicqdfSeP0kLrQonOTng4GAu94yr47urHX1fxSlr68vUQggTqJshHrkZsNWGc7dmD9ek77yg
2oPezPO9TqybB87I9ODu/TO/6csjuvVoV2QyeiWhyy/6nKYrbS9vDnlRGtBVejSAtjySvFDVkFYE
24N9Wj9apnLgJRcqM8gYpUjXMt6UNBUHSVZdzJsUjgmoE3hsUDSef3VRCkW4eNuIuZU/DYN21+Cn
SKP8biKUkuPnLK4U0WQsNQe9jMu4pyOBAaHO5fFoBqVXMSpGV9rzApAa+D5a65JPEesRsf92GDMk
7mkMcKKY2hS4hhARSzXnKbxN73rCLr6n2Cn0u6j1n9qD6WhWfldwbb5jNx49SdMi7vqsLEGLllXO
cfswULGDaflZFs41ml4W/AoJfAH3hwezbmxWqp/jUDtx6lf+wO2QiZ1AMsaWDElB64LwnjKyMETp
L2051WRUlwo8RRLrafHxI96LmoZVrlUoJM9Hicc4czz0QlvXt3IhCw34TlNEui0QxTv3dHMm8bad
+ywR/RtZTyzvmxqp9Yv/JKPxVfYzoEDUcCGZzbl1mDc09s9qHIvPZkP3WBVjlC/kdbL0t0Ewvn/c
wDgZqvSYUuCkKkVsBnA0thdFIsWWCyOZsxLPO0MLPNz/d1v0ugCEGvbStcuiAP/1N+zfgpQx6xBH
H8kSv0rsCf4to2RFs3FkSs2R5M/Mj1++sjVMXIYiq0iYwxXy43MRUZVobe7/TG0Y4zjkDse54EDA
JSWbKUmkRRTg/FVY1x+FjjXVm2hnaatCPZnvag0f2R2F7Sqei5IPF2AdzwKdPobLqnjU/OAouAzs
2zM3olT4jIbdMEmYFi08V/+P6wDDyYrqemE9RdvZdGLTarhNtAHkkvp24qHtWxTaAWMZTmKdTbK4
AdTEi9UQdtJNCb4uY7ehKAGXhjBtxr1KI6p0KHXigWjwefaNGQsDWRRYQwTwCEjWC1fZnCdG2nDh
1yRuY/YMn9L65doC0W0LY8FB6GHi9PmKCWw1k2DRpgLllMHaFfZ06ZCs9ijSIt6wM0US3orPTcUx
7Pl4Ymza+1B1Q+rg8s5GfULFaHDIDCCR6nuCKo5/OFb7kWDLxMgn0tQRWtp78U4mgtE9P1P8WHMu
RMKWXqV5a/3+lzAA+4SUOgFAfAZpIfGPWikqw3Gf2uSMy2vUYljyei4tHOQGW69TOBSxaPbuqkuG
eNfY1HUnZQZLpJIfu254f7EiOf8TKrRZZHYuzcRt3ponO7oZFHgt1+nVVpWueQhgR3sV+0J3qTuf
P1CfUn8JzYuMhuhSqSpFHvM/GIOmVd7wlskWd/ilH4G4tR/8Bm9kVgBlzLXEpqgk69JrONKNvXfK
qZZmqqCm2vjqa57Oyg7Q7grYWA3yBjxYc7h4DyKlH09wCq8Iwi83j+hEZA1sD7Kbts50pkdcaLMd
hNdMELX9ZrLI5Ji7lh94ha8z1G4VaDuKu9N9xMMbhBMhmMWe76SQLwn8wEYGlw11Qe9m3V9B4ZZ3
EEDfN7Na0fqIqzS5uGBOnMvvgNb6mpnFZehPKmqszLkBywitvCDfT4/CKMjGZSk16mkTY71gJd/j
SzT5ohtMXV1nM3UVZhKGgoN6FvwYrna6x/eMYuhKvmeC20tuaf4yFA1O7yc+fXEPJbdUG6wvCk0J
hOjuacR+t5gfDlFRELHTWbambGTnfWcsy+zi7n7sNWChkt2lB3VL4mTEr2Ucl6LrtyjMsES6JNPZ
RaFyujkyXXEOGRRdP9PjtckuLmAyistZXTc2gNiE4w8xfMTW1T3XeyQQxu9RJuxP0tzzy4qx8J93
myOoBfSIBPwoxuCG8WJQUmOPCaorDzUVsAAu7auWkqbJdVMYLrb6NzV/05kgEapfRb267rVcgU/W
oI81su7vGP01BpRdv8LApbFKDHvCT5T0Y3jJOB6km1oriGPIP+wvkPdJ71BzWXCV5jq/5BHSYVjG
2LDT6ViK+8DOkwAHxuAdHJlqOBbM0mQoqvOl2Qux4XPNwv8EjCrQ8E56LTgeU+d5l+bhWaTeE5zu
J/C2RUG7LrfaqrR6nPdyu1tQYezD1bxz3xuYniqNaSiTeB4ul+6E/npy1Dj7FOOyaJXppApa+pRG
hF4xFX4+8oBI4AgngD59asA2xVSYHGfmz9GlP+SRQbL7sA+gBpxtAE7LuP28pLYffM/9yhCTsqAt
idkTMy0yuEeZurBQtxVvEEFHTsHfcG1bM0+IzYulYLEdAZ2PpmsDgu7/VKFzg6LBDVhz1jGspG/D
qNQt++0OCnK2CCN+9rJY0wzYaCqy5c2NuP/Gb+iPtypUwzOV98mg3zYJ6qGGAWWh4SY3UJXbFDVW
DAr16OnUTZmLYxBWfDwWsb3jUbO+foNld1d1f4/5zS1EDp31g1QbOBgiBcae/S2VR9wcfXViDBGS
VIRBhVCMkX4wuOKQOZT0sqBNjFLIz0G6ksdG+lPHy0ZNR+u/aJEWIf8QZTPju9j5sjmKLnqj7Prc
HNxPh0hQBn3pzVbI2X9UH3xuHZo5ALDpumMg5gD37+gidaS1YoQucrBQWaQ1KxV3NKb7w6OlME1T
cNI0YQOxzOMlPAKXEC0UQ5ky6eX/TgYJ9NzHrrkG/tM9BhPeElNYEWZ0tXFUuoT2pwzvPuKt0bkc
1yGnRaeUotHdDiJvQ8a4gEclJaFKvDq17E+O3VTpUd5SbrUfVUpguzWlfxMOQ26PhAawOuyXi1SO
uTWkXnkzFlYZpmxg+JtnRMxxYVrSkEsTsKBE8so/rWRLLJB914KAqmNHcqQrSBhvxhT3JrVgX7JK
c1ROeoYlGuldwlIFTeKfXOJU5Al3kZGTSYtPQsF085mhVN2gufzilq+KV8Dw3N+Zk+Tm9mBcY8uP
bmK+v9BRaT7Pkm27tkRK+HhdjKYf0AwsfjBtisi1/T/nTkfoGpKJTVSVCSajRDjrupiSmIxENcbn
36HpXnq1hqUiNRcgagfSg0CD1LjGRrNIJrNw9RZJO3sl8Xmy0zIyXYWJIOvnVp/HxRfbqoq8iMnO
3tL7iDBAfAKzbO+6maEQmgewhJWNS9e2DNbCpJqlIABYKUiMxjQubYvufHIm7A1EceLBS9gFIGeF
nZiZvKYmC/P2YfVhcmoPDYBoP3L/1+EHLW2icLfi2YQ95c2HT7c8a/xOZeFdnNkMsgb8P4NObq0P
DuD+YqzgieAs5EdNngLzh4MuIajivqPqIuBh7Nybb+WBaRilS8tI6aM2n1xWykkNwj4LlhAVcWO1
yYCTii1vzyfNDtqMtHTUmY8ZTCg9na106PledXysw7YnqxrlIAwRKL+BlWoXJq2vmoJKUP7ViE6l
tcKwMma/OjDaRERNjmqPMqwoT9arGwV8hB5KZUahs9PwJ/7Acsn2cVW46/BKGiHieojr67G56eVe
r3wvi8vwHjm/Wr73PrBZNL7MUGqsQEZO7wBtL1jwq3APguXGuRcZWkkSWG3Rk4tZN7nSqbw9dL2+
bdctLWyGoef7tv1bgIh852YXdeZtDc37zrUvMJmQ/qWwy1FEDLjsD2g4VcuavEJ3Pi6OSTuKhOxT
7MgCaKrfhPsjuexypdMjCwm9jpj9meptTod48f2ZJDMT5BU/Gs0vIsT0eWFQVBqNoaOAv8637Q2s
6PXW3zU7kLkdDJNiTbCaf5qcRjkWC0VHN6eoFeviyImL6X6mYeEw422iMgX2frai1KoUNKI45SoS
5zmCV9559e9GM9K2FkfSMVnx6v5eVxS+94umzx5+3jcTAg6qpFssuadWxcsCBrBfVFiNbgUkPUSE
1ONhNpQlnYCXcOtF8YWOp13SgJNOO5lfRU2HHWT4WjREKQzmORqcX48X7YJWxuqFzhsWqHbW9xT8
tSVQFIVyP/f4EZvZQL+TIECa69WCsDoAz0lh1eXXR+FlQ+NHvK6vE1gb8i1JO0c1hrLF1KiFE8bE
TM4kk7ZKA8sYwGPgX5SIeLY2uDl1uIfQZEEdxycoeUUDZvn8ny8afrvQkmoUTIGoMj/yF/Oc/2gh
RqX9ENShYMSjHyP83m4jDmwU+P1d1TIzKFoasOokeMQsxTCa3hDXVthMp+z3k6nxhMORA7VWC7Uo
Y1FTGSLSkfB3NMYHAzXi5cTjhDjh1uh2Yn89qsSggRL0zm3sDAiBIooZdm95uEMLBwMyIXKn5A0o
/TwyedNgyT7CofXQWZ3M+oikhM+eXlLEpq1S8oIK2oo8UJgaYINaKnzXeMYGs5FX/lPbe6ma1+Yz
UGSJzXMkzFjfaPkTue2murthTJYtSvvqkN4sv2SRKZDaosG/lJolrySBrCG3vjJYrIbEzaDtDIM+
k9axPN79G9qabREmvssBAPvtxBDW/P02ewwoQ+GPY2KeDlCuULit6iTdPZVf1jRsifuBwUnrv4sX
9GBzgt0Idjo6c3Jfv0ew2+gWNfg+KAoB++vYZOyvcyNi25PmwPsGcj5aSBB7rLB6nYMebdT3fbGv
jwENhtyVjcLiv1Hz3nF9WeOpciNUK0RSRit9GfbYmcH6ygISflaAiZLT5TyXYHELkZf+1CU3tpun
b3MNZIT/hXeNS4ANpis+uDa3NJ03df9LUMrKDskM/ne8lM34USPmf12wnCdHW2iFeJA7sirX3eks
UbEB1MX/+oZBAodMiEj/CJZNKAbIjdvRmoz7Je87/x/qaQgAWKwLLjhjpK28W0EyBe5leZkgG8ag
p78Q0ngwLYT2boT9W34Tt03wopy0dXsQm+sqNzCI+BY2nO0LIIJc5OHnIl8RelVHtEENRZ50OQm7
K/Oqc83w3mMgZTOhdLomvRXaw0s+IKgtoGgKqcIrpv4LfsA/NvigfreRc7NEJ0amjTSsAgeXapau
t4Jydnj3x+e2r7tugCSstQ4r8YrkRpbsmp3AQs+DeEZyNYFi/lv59LU6Sf8QlLfnROANwJPnnef4
eRDWVj2DO4oN/3gAjrWSpvRmYMTCuuGfhbwVAmcWu/4mx2OxFF3o3xXmbQOg+NVgdahY+PD9iHgl
LVvKteWcnZHBJiHr5I9WZpZ7FTZJ6kMTSeqSFIKXlN0jT3Jxipb/QNOXlZLirDZ/9uAIw3SB7x8R
0/jNPYryufqCy75LwFeiPaL+ihZj0HJQ5cgSSQ/H3d9vDO1H4exxr3IzHl5faqCJe8u/2mRIhGIT
4ao8y7bx69WfePoQ4mPDXbOnLGYLI4hutThw5Rf3PdTYgL00QDvRc8t/iBAfUjn3a6iOzsV40mWF
2yPiWSh3Lo2Zw83/skKfWfp/+2NxYENw0K97d4qZrjcJEzn5sBxmSDuPaKtnF9n99AMfGLvTXD88
sx2DwHlTyvpqPSSZ0eIyOCqdPloGXhQKaIdq7HTrXDhpMQNB+axyyF6plKAzoonOcz6nSerVaCfh
CXSqFyqyyyCoKiNAxl+ls2pBpA+bWza4nOSEG+O4rPK4jZFYNFKsV64d3s1Fuy3+FAE8qCQzHYc0
+kI/H/9dugeUojqDYs4OQtvH3UIiYqsCivzB5+wdjzJawswgLfSuaV6q9Mw4t7dF4pHaq+9VOLEK
hYZTXoumb6/LvqwZzaMkl+idmbnSSl2sYdHyv5RMHz94b6lFxX+IvF/tG15kXwQEKn2Knv9zxqBB
flyrRJNVnqjwNlVyfKsg5UDdLFsJCInJ7RxrP0nKUZVdaHe35poWW1M6vn6aNdh9pBFtSPMO9dUN
m983QF8ZPfs5FHIoKNsD7SKcu5kKFuCsRn1ybwKYrZk0B3A/ShGPHKPdI7cEmANello9owO6fWFR
jzwXspGGEAhHWS6fuK0d4cjh2uQTSv0Av6ztGxsPw0c+TAsSQvx9kII1jzOhYTul1uYP+twdNkTN
dVLEyczh1MBW9VQqheKn8tLzn7dfelgPOMfe2Tm+c7LYkALFlMJCkNohfNMMmqwycGQy4ewHvqOO
6Ek3YedFG+tzATciHynuFtlc6elvCybUNSYrvRsA/nPQpHPz7YNSaa3uD7dRX15xfQXBsKKp+izL
PHK2oA55gaKPkP1ZzLHvPjr87CS3Nof5pPZO7+70U99qlIxka+TePFxI8bC9kqpNUkhZ5sCaXzLT
JIXhHB7eyget+NoVlH4+EBKYlK89m3Ml+9htXMkPhGquRcnxPrYEfXW/3i9XTjHouk4uLLtmusib
yUx4kKlRbMmBSizkRu9+sK2XaSpww6/WlsXsyEnAf2E0ncvf7pJgbMB8p4P5yQPg00NQXW2CLYWZ
r1gslRLvUAm2dumYH6JMEIhir9W8QUcVRWBF7sBHcJc5/llS6P4VwB33l4+61ap1e6vjM4PV3duR
QmuSYsD3spGS/leWhBe9XWL3pwxovVyzte1KuBwSg57GD02IUjPRbQMzcEqYr2T0GYzUhxoid1AL
7q7oNBl9+N61Z4FZPciwInV+6kwOVvVYem0ZU3iG+qRb+kHFAajv254nQ8zzATpuO/dibmPPcEqV
j7Vo8yBfWmpXEcZOFrcJgfqfVxjNGokzFmf2Jfr2T6A81ox9KJF8R0Q1RKT/xuPwau3jm9/ldrCQ
IdGCFyvjd1tSaVlS5mC35cqt5ot47oGM3VhJFBIwt885ZXsbhoh5UQ61vlfmQmBUF0KkpcSObk6h
X0gX+ws4lpFtcPeDoYdhNI0on/pa0dQk7RmPeN6va/+HPs78tM1RjwH9CT3qGmPvipk7w37Cxb4r
swrzGXiRJ03Rc8JWN5VJ5IxkSt3L/P7rpahKxC+kM+bCybO06dSeeHtXKbLxrBojzDSjUHcWMmVB
Ej6Qkj319DV2WLc8xAZamedsWW5klbBIxnS0qhoKG5ISd5q7o6bj7H4uai43zb+zzfYSx8+QOYtX
7V0ZVY71zL7YfHlrGK8lkVVTzFtTtmghVFkUzFZmhXGKCIclnoLf03fhPhdmo+bmJrUiDlSJIOBi
KI1O+AQv2Kuxjo0A6Da46Y5grB0ev9rMadNMB9NjEJSgnTnPhQEIP7imo+xmXX19VDASUXboUi6j
oqPB9AWznIW8gXT0qa1K4m3o7Jc10qMeX9zflsejAPrv53dU01aLDlKOg7ORZFITQuwCq4NisvH+
XZRt6L/EgYqWTulWRfbgeSv7uKav2LEebbztFMgAx1FejEFq9Q0qDp1tU3qMqH7x9HNq4IC6tWPl
Gedl2/sqkr7i9BiQLQXrg227UEGYeiNOA39DaqCqh6L5qWJ1jn5QVX/qQ9UIeEpo1A40wq7peegw
mhVlxxA0i7zESoAARlIM7bJiSekzYjRSf7cdbyllEj4SXekW+2nR/961h9EqgA6FEKVHAH9W7jrh
n7UTfpWUiBdbazvD19bFJtb1cug7AfgRp9W6PXV7WNpw+86MFvoliX2Lhf2ivTLGq902GQmqYldU
Ebl+if45+vCuKMUa5NJ/DLlwz5TJdR3/gp9CFtcLwCnoalkHie7mq7r+TcpUgnHWxQ8lL1fs3H9N
+7KpOyO3/QzyPTZjhtRQc9X0BODHYb0Pa/u4NORYTV9o/6acvUbQ9kKQMn1+Pb7YdSnmA9jFsDlL
t7mAdOwQU0oo3XItcxgYQoCMIo3UcLHGqGWU6bIaE3J4oBpjkOe/jHocEnPePuP0wKSp90gvYKop
Po7tJyGqQnkkceeJtUm65oSLxPGAwsW3Hjv2FAxGvattPWku2oPlc9Be/tWcdbFHDB6Zp5oTGIwD
7XkTHIfxlVCCA5FVw+tJcvCx5hXAOgbBBYgh4Jv54dQfOG7OvtDR8jSaVRkCEI3Hw4nazdeT/iQb
R7z+pDJDe7zfp4/Je1irBq1JVtStRTBM4y11XfZ9h/kt4BGIenkPZFf5xr5kAN3nJIQcNYS4//yN
H+YXuFnMAHJUwenoXHQL+LldOXksHYhF8mg6ACkqxHjrBtb5zvXVO9XXEa3MNWRFHAEPQNm4kNVF
oPGFYDR7vyHKd3HJoBDEe/8tfCxPlu1mMdyzkAqAbTx5SBpQu7qzEp1UUMfSCtvARNI8knKbpoNG
F5QWxUsqwM1Xd49PEPejuFGqcym8mFn8GsCIBvDw1BfDXJtPItdgEaxwLgksS20N8CY8JS0bbPA7
is7XabfkbP48AJeOx0W2LYjdoPqChrRDpVl1EXMWwhVbvIk3GsAwKYR0LZOfHtq9wU4Mp4KU+0rQ
8PQk6Pp3L8gRH26HGm094IMqlqD10olv5NUAcfZyqdelGA6N3cha3Yfx0OGEiD1D82eaSNAcE8+v
tCvPpxXHMiEOwcK4o4GemXdohmtceBaQ9DjSlf6lRq8Ag/fo1MQzLSoTPx/jfAFBPffXTvaqxsgp
KMFhcyIjqMafLUyikqCQy0SZvBMOhN2dt8eCoGIIpNI9zJ54YgiVoZ6qEQATn1hoQxtLBMZ62GpY
YU4WrL58nMRNPBebbHYvGJiT7ni8dJGlgaJvdV2KbM/RAhhT1RzCQHth/DVHxLsaSqLgQmYMFAIH
FjMwALVja+Zc1BP8s8W6bGzquKqw7u/ieUimpzJYgAJ8vbOIJzP0EJTkXBij/fSZtJy2+bngYcIs
FnaB+Ov61R9T0mo9LXSRbP/hBZaScBrtA7Ng9VRBiS1I946S+1GmZD5jZ90p3JVsMvDHsvkvIvb3
VEjVKfeebcbaBpvgdyDQxNQrArcxUqChjvuF0vp+fPyyt72BCKtNMgxLopvqq/VNHhiR0SlM5U9P
9QLNIgqauOyTAczemqZ6Skocj7d7klLSswidjxAIkgcOB61W+yrmZhbeR7j47frEBKXsjzfFSDv1
DoACF687GjV+4c54oipzS2zNMih8iEB0dvkWmK8Hnim8Bss5j1qxfVVSeehJhGIAQ1YL09CnRIvk
Tg9fJ7mZl/qZPcevLSNI+QxAilyXvZR8u3paYzy8G6O/3HqHMf9Uc0MGgeEtePGc/uhfYgZXn1ih
oCM3W8x9RvyonR+TH6LkKHx514nnAlXgdtJ8Fpky2x7z5VU4yhdgkGKj/klbKybKMa7M5vIkwchf
RQPUBH2G4IBGDw90Hh9wjU6UmmH3+GtTa39Q6vHW9GWfSHhCeCdi68/zpyjQraEZdc3s/t7Zl6Xn
tITefCu/RSmRm/x5Py4UcNOBlk3ibjC4MQaV4Y2gljBFK/lIDgE/xi5fWZY2a+JrF2mVLCC/TAOv
smon+rSXHUQDHeVLhWT4kNpcMQfhVfS21smEX3hPYq1l9L1sfW9mi9n2UK0xpAcP0jL1U8YGPiLB
KrpgTNXTybds+kPL/KpOpdFGD8pKART47BcCCWde+PDowCoHiohAU3FEgkdcnG/bF4iie11n7a4B
073TGPt34YR7rBxOt0WA+HBvqco5wl4yimHg4zCCD+nFaIOEexZcM5ZQCwYI5O3NY+K9uTh3vkDR
19GPr0K/y7mqo/ONMl90uhLu5f6gOMeWKfiNlKw2eMaFgGtKBkz3SuQ1xi3GghvLSqJQfUpYYrnC
dMNF0Fcr3M8lS7GugdWSM0tFZoHDvO8EUTab4p5HtyaUedby47sDKLo0WdFXW10130AEXh2hDaD8
E/xuijDCcPsSs/1H9Rw4dYgbHNL3sxKO0KQjVwCpp8yX+x8C6f8GbtDUxHlSEM1REJbfubXoBFHC
QCNUkZ6uF3CCuNGnI8/ZpG1plm+lu9zgEUtR/OT6U/4hl3UzUSQ+c1R23taSAZi+Hjruy7JIG1OY
8hVjB3RgRl/c4eyGBzUyKJDkNkA+/EWcG8KIHrz7Tl6aBUKTAaS0Gbxz0gYHS07/w9KUKTxtPZOv
P7zhQDqSGtS9/vYbkt7KSfiD23V+H497grPCBqYKUnnLNgVDd4FDbKZBQIrsUCPBe4QSpVpnMJQF
uXyIJFT/z/2JA4qDjM8UHUePl2l/kDxGZv7kwl2q5zBDRevd95LrEvfCz/2dEjzfsi22RBZwFECz
rtclPyqUDd83EAU25o8F7+bw4ArP4be+gQhY+Qhj03G18s7yWSC8K2rTByCXvWdZKc9dQA4N0w0u
indQzzQAo1gSQC3xzuYalz2f93uKvQt2tp5PWfJehlm6xiauf6kVTc9coCzoeLoopjGhYkCTUJwX
Z9oXoEAtlg2ph4T5xlVPov/9GQuGFMjPVSmBV+T4LFGGiFYcu21jyYgayWIfaSzW9s8XzcKG0Cw7
Cv6yg+dfKx3NU6Fe4FfQJd+VY8pqjLm4Tvr1EqlRkz01AKMbkxdDsgJNy3jRcfQEMjAUXziXgHV6
c1mZApukFF+OmG5izAaL3Qom30MBdns+LHzJ2ZKz6B1bp1n/sNDf8C9dc98YMuhSedAlaFxVoH0W
tjMeRnAFqk2z8N17DSc59N0jAf1VhrcuJw+px5Y0EBnYxNuFAZOq8c2QI49pC+FdNV6iziZO3uad
38udSe0hu1pjA3urqaeeyhKuNS0pTKBvW266cWDROxcBA1hSfvVzN1lAmh+l/tW23ZS2METdgYlu
C8YepvvrM89OvoXb/iYfo5WH1G+uBAjplgHKpTkvG5cesY02e6DE2XHHnaIwth5xJ9rrKwx7bxDz
yS3UMotZO+4GXrwKJHpWXGc+KmO5VArBAeT7o0frL5ClJtXi0gFKYmBLmy5Ki8HJn08ovyxz3ge/
qMzacKNyjuHWQmHK9EvqB+6FpCXX+zwuPqrXzx1hxf1ENQtIky5rHLanIBXiHiPK08HHu09PZ+hG
5hwPAzvdsbUm/6NXsKYC7Nu827RJXFCUfSycGppcDR9lYVr6nZ+jph4nEuIrDqNJiv1KkIP2oKfJ
sxXma3ZZNWO5tAQMycMlE52bdPJJ9EYNpwQEko8D/matD51ocqRigRXsbiHj8x8wpbJg37Wg7D+G
do5INwwe4m4pLYGbawr0NuhjJochwV7QskqhroLNsEeSUTbIm3HfwBVFbfzUgUtojzk999CZOA+9
dnKIUU/uI4OHFX6zOtDGHSuAjJ/fQVJG0vwZcruyqh6QKVf1o1hodsWS97ycMjK4hujEcbvmKxyn
VxIlnT8XbUb2dDcdTpy2FslbIVA3Ah9FV2VPunghzVlPMrwCJ0Z/usQjqtXFN4/G3Vvw3NvNW/bc
z5KPM+xDHpxMYX/WUmua+q1/9eZ0OPCscfXXJDKcwmCsonhO5aaG0nmbAJqisLu29offSme+NG3e
iIJDkRWaWaZWH+snNHPRJeBjJhYZ00msCFOpfQ2OKDEI9qp9z2SYPKaQFL6hY1VgvggmnTTxnCZl
1/XONPIyJvQ0JCmNXM/g5NCvzFgGhXjuw6FXs9N8FLmgB5HBozdTMTNI1P7s0WbsZjzYFltFpQx5
bid3t6bQorEFDMEoiXmYl8ib72psMaQHs7ibaAlmcrfSlZYuA8c8Hz8akS+5pBHQlltzJyzYDix9
aCAkpsdJoqFqQNKRArnaXQlhTJtE3U304gI6PWQPcMrnuOZumHfAPpnFIfBpKY+oSu5oD6El3UH1
9j4MuBTGJdnjixsENBunWMpktgGrRDmckOwni7cBzNMMnNAc/mXoFbuFVf/S7QZlS6pTwyyzj0O0
/UYLRBzxAvEbqKQNsAM1ZIEwziSmZAFMAA2FuavtNOPq/SQFIfWPV5xKzUzzOtbKJofFyzLkFAhe
g+q09r2gCEFJcWDcLehn2OBztvv6aEAfY8izHa3iWrH0jjdL4fgvyBztGEgqjgF5X9GfB2zNRJv3
UQYdcHHXo18JjiCVEAztkWBFFKg+1T7Jhn9ZBOQ+5XebmNSCw2zwaucRMgpJ7q7fubUOFqBcBaQK
oeRNQ6RtlveQjpxYZn/XYSzXb+DIcSmKJaXdVIP3qLKblSnBEY+D6auzDmxymM9CITeCVot2YVZc
V/sBmNzwuwdirA/ZUIMz4GncAZLFN139tWRiDvQ4OvQEzT06rHlV9D9TY82riLHnpAn0YImtTYKj
D1DdvjSq3rUABDfWp0WrTFwDrQXTlUdh7+uM0GVcSHpwfCNmSH+ZGxs7/iCSRaWjmqwRJGl957Ii
Sh7Dwr6XxKMAP8gPep5x2sLVhX6D7oX5QheuFNTGSzOg1GToDdKCATEZvGyxkQcV+sa2YVi34jLg
FllsGCV5nNDBv3L+59mEFEF+V1wmdzN0Ma8ibNdURwuGTQK3kKIudY0jCuMPLnlrnwDsDKku3L6/
RjeqNmtyE3rSiEYeIulrt+MqV6CZw8rfgtAq4YV+Hr2QO4XpeTW3kIAIOcxf9Gdd4bP7b4Ke8h1t
J5RawUnL8E4z+8Zln3AklO1m3m3+RWwV8mE2iaHu/ju+QSqo8V+KGcD6KWj1eESE8IuHeFk+Kfs1
BTuPX/xlOgQcsAJts/XULHRv417Gs4gMXKz8zUIqj/2D4/LUm354myQovb4yCGXXccHyXmVqnNJm
ILbJTZ7r4N9dilR4EMU8Ej0Fl4rzCvdsJtJ99MC1J5mLz+tXyVxzrYWNXnRFtRhtYMMtqpJT6qRP
/pMATlLKDqPBB8AGjo4mTP0daGBtYMxVEOB/sJL/1SnCF2AOneZ8EZF2pMoFT+Qik6SIhpnVYJoN
57YF81fFlQHTpP1n2UquQvVowsaRwgiBriRSPC7BUSwLF8htQQklDwteb1zE2cWD/Y2rhn5G8+hc
d6o/CPDlA7i1sxMsG2BRn33zd2x4VfgQn2TX9nJPzWFzDBzzuBzfQzDbAXEaVmHianRKq1P31dkY
1HQJm7mxsj1uUDY+YmAMTg3AC4TCHYVZiea/KD/INOaRQ6gOzEVUPDABra8nbLzpx4kehn0eOVtX
tkZ9Mlh9gGI6gGRp+MqYa/M/JDqsWIkLHt8rjfWP3n/qZbDYwNimiT4MAb9FT4k6siwUUZgpJXbY
acYrlJ+Xf/dJ7bzPuBGgW9RSi2Dtz45Lcu5gr5PQ8St+FL0IaB0E2zQAtoJecTMznxAqX8mWNp1E
cehWI6sHD1wVPhWX39GVAOz8JBFZf3vSgVsfMgKyro5j692svr4+k2DncgdG8/PzIW+a/M4YkY54
+aIdrvATDXoGe6gTl9A/09WGe3jU5v11Ol0oHfzhXrom3KYDDb8eNsW19Vx15eifWAGOT/mME8yz
wDqehPu9Gq7QUA6XIplH8Z7le/6f8Z3KvX0xUjfol1UOXIU0vjlmPpDAasydVuovSfNdYRygkOKH
AQ3QSgb9O0hG1DRh2DEVd2wX/gdrqKih663t7FtAPifTrtHHqDHeU1eoM8G5rKeOX6kOhJKE9uFN
gzLy/N2KFCjiPvJpczfFWnQUAeiQATjEZ4tpeBKtIW8i1osqnQ+uVbWwOLRS+68etFEPTjD5Vy2j
cCwYhCdaGgKorq2hr7lstnpAmqGKj1njeZNukDx7IeFwALe3UgXIAq86gTy5z+VxsH+zLwSE85Jj
Akk5f4h+GrjmCIDtQm8XV9Ml/fVRaOQA2EvZRvA3kZOvg0u6HtucrXFzQgnlsnCWsDYwNK+9Zk/9
SPJ9IRtQafM5T+3GN45MiYCFRK163owtift8Oj57tmjq8fspguPUrWKsJm074F3RKTPuFudFUniw
557QarSv2+rwPS3Bs7vpWcogdJHFvRYLLOygEboS8AouaVdBcgtxNi7ZHClw0YQOsZyT+xYC0c01
N5DNCwdstPUctU/OtZvD0RSzXfCmf4hqr17djA43mGPwlBpq52HOiorvxlCml8zfSC5jGiEVpsvh
BX7wELWF/1/B2HOD+p0Wtwybz+/8U9DG7grdmaKzMczNyi4li+QkTQhv/AMJpJrlxzkt0CoLJk9v
Lt8ZMEB+FApxQCNkn2CvC0NdG34XaXgqGRNRBfswj3mpREmvr7nYC6kmt2/nhFN5mSWNWbsfZsXW
nNBveneTC9lat/tDGK15gtht8SPQQ/AUuPTO/LZu0ME/MhN5QoDcUK4vpF4Iv/VxlFmu6AXA0OSt
jrnr1TJsfpQ61SaW3ndoWsCitiKOp3+ExtDZT6c8ikXyr/HLQkMD0eIsWiTslNPi0SpBzuweWRFr
AyJxI++sQvdW8c/ZnQJEwoL+NlLq+Uii/4lR9fuGVa8dZ8MZBNEe2xNFcfJlQ5ofCu4g2iwXyyEx
IOoaPyhsxYgMduQflj0fBIVDaTQKqvaE2IwYcIsRYeUoecYrYjkRVLrViuHTUyQ/Qx4geYgjtJQ1
p4RlaWjADTnQdpSuCwZGytIbRIMrc295sBUkYVcyC8/spvNiO4E89iQa/NOZH3E1FB4MBeMPsTE8
RD0jtsFRhdapzxxEtQgX5f/WW1fHaBhgeA3XgdexRVf/2KOJ6YHCVWpz9fsE3zdQDBVUnzW60NC7
rpwrfp+fGjC/q6OXzqbEi33Z8s3sbvyWWxJQkuQFWchHSm5Osm4yli5LHM8IKieeqQzqwBFg8UX/
tzO+3a/C2jr32qk5KiWN787z+65qr11K+A8/EFf9A080ZCVWP14vjvrQm2aFn3vyyqPuTdd4mNgn
GTAJeWF6SnB3JWPxYFmkQf2RchFjKySUpbeeYXPZ0EiK6IEy7Qj2fqAaHdU37WXcAC8+7XfWDUL0
6nP5dTeFZ5fvVhT5/iIopMrL+uUUmVHq8nlk+w+5/Emjo+iml/8W1SswHknPxqnIweUPYHFvKEXR
w4hqaKSFBWzRpfZ2Z/G+khXh8ZyfAgU7YEWF/UfCWRLtDYDagGJd68Ss6/xDuN2HNjlMxQpvaiSt
rRtvz4x6XnsqMlIhXSNtLbTcLcs1RwrwdOLoFA6R1TZK4a66/wX99+6xK/Bb/56U9Kl4OgyENVFB
L/RIsVmDLfuRkiqK2nMbgL+HRCJaZhCptDgk1yLjyw4rjlOdg8RS0aepG+KU5H3A6Jc7kGfxs5TK
jdIOTvY4Zpy4PWeZluxcCqE5XU8UWqisjc7F+AOaVK4VEQZi1UyhUzGQW4rTc4QDhIy5sL5luez6
NMPO+Z72baszT5LcRsPRXBgVWE/n9AWgvHKe3CrPOIfSccVUXUB0ONcsP/Q/RhZ7z9a7fwwhpXcl
SAHYmN8Nw+GcxMkh0GCLSMKPIQ1CqHbwhAOhncwvCLRyr0GSlp8IrQr6FyhYpkBmln7XCi0qf5su
boBOg/D4oJCtls122wLSIT2Se3HrhGoFkK6CvQEFSSD5HGwg7Clbjcfq7GRdtB74yIhO1eyQElw8
knBnFBKnfvUkUNsDz6u9QOw0G0vy1madxtn1gF3domW825Q62hleqg1x8R5nD/r8jBu7tognAreL
Cy4ihlUsKioLzSxMcMhJebHssgX+UMEAiokrA1cw2dLvM1T/FAZKVzTfphfbKlK82nTd77uHQ+pX
y5ckjCD6OnUr1kTlkyM027B5hMxtTPUBxCRpP7SVuNaf5TcjhmA9ariWQ3Ti5sN9UJKF28OsPaRc
FGvymZOPQ/R6y9FMSw+7ayI7kz0ZmE7l+yMKsqgVvAQBVglhuVHE3v0+GxxfM3MaU6HuI9yxF+W9
dgUhujvl5fIsSHRM6Mt9oeIGUQr52CevnBqzA2Vb3RqZhlMXfYqFNMKi8wALWdJyTQoiuvqsv1F3
TJdUrOB/8wxFJ1tTt6tSpKYL2NFwdqokZ+J3RPPvfC52wO9+SCRM42l0Ih3V7Itkzs92B/zBTeQP
TNb9aTwfgRWBokmTr6Io0lPsIvUW1WclYkn2wcCG7NobnlB2vlOWhuGD3KI02Ijqap4Eztz6fslj
QHc+lmSG01CiKmBiWICYXLD629QIOMBtG7JarAmu3c+SenyMTrAXp+6kvzD9DPWhxSH+oJOa8Vkj
DMGqrLGjIqukFxDi6FghDIdcDS5CCm0SeTCIkI3odI1x/cpYJHJT8FyEdd3w/OydBChqKTAMb8Eb
Q+b03M/7LFzdFJ0+oQNjz13YBU6Tqyw6kwKQNVMuJjQaL1ixJ739QUHuPcAM58T+gnwHZvIXyuK7
7icbNFioYs0oK3AofV0eZV6vOTe3+UTKnqjMOFCWZp+z5LWFGF8vcGpb340nSYRi0giCC2ZHj+KJ
9jJFLFEKhKzjj6JMDyz8Y1/WGh59mu4HwEwzYCjSFmQxJYsAqhb9KYNhJqKKhzrF0jxvvNxGvxb8
2LDNTSY0r3zrr4Cha0naaRq10HzqsMiR4BfzsYOadVaJ9BVQFuLM7pxM+XTCQnLLbmMBqfJfS03C
F/4qcKptAFotn8SZonDgTydJEa0/RHTx8H9EkoWZHC2RNfj4GyWON+FacyBk1j0HYmUpKMQBUUIl
U1bHPcZKBJYuSO9q2Vb7qN2tEHMd7N7x3ueI5gORlB8cWtNMCZ1D+P/ECkz9phtgQQ7csc77gnWu
cY3D3CF6GQoGidJCbr2bcLtTCJTZj18hheopwp92RQsjRnuGogOpQQOasvYcruFD4VjCQ3BuB/rX
oaK3FXPml8ChB0shHbJteiQZhfByvP9yHZVRNoHsQfKa2HYc0vTMZt+B1HUL1UZS36VFJCUN5npy
SpW69SXTUoJ68udyTDmTnMPF/qsUjiDyZnuVIR8qJJh8QXHeew0D8LKBT5tU2ORhgd2+t9sz7Yxg
VJBtfYs+7YsjES4OoxY3zvUUS7jGfwXTgul5BJrYrWeGCbIhOasmwnbXwVpBsFi3zp4mAnv4sQAg
hU8F/AL7HipJQxHJYLWwIwoQ7v0WgZbwmq+Icco1pvFvnm+BkzG+7BTUp/MYHr/oPJj3YtHSfPTi
8CtmTLMGXqEqYqiCkfDMbIZVLYC+wAF1vK+R8rN8AonOAvj7B3eCvBXaj5IPoAD1ceq42XL6R7Ef
zY2MNVX8+JoAh8Jb1SsRcRLwmSx/KPMUZYTCyT1YujGHdYkIRItNT4Rs2y7QcoNIPhik9k0NhqBN
xIe4gknhh0rHiLFw7GUhl+8uJoTu6PUhYaLTcX0PeooE1V0NqYig5oRcfY+Qomhvux7+BNQ2uDQQ
9G/1mO40xZoeLUZSs4W/CLrEiGEF3vtFmxA5UnztWfiJ+/NZmhrYOVgxnUWXlvlhc3vnI5k/3raN
Dji1+0V5GcM2u5aW2zJHHwxMQjdkOH/kMOi7vcTNrHxOYh1MCBQjIRkSWFek4I+mmgZrnOEgU1nc
pcvqUEnk+j0/HsjUpm2+kPMvn+6lzZmBFVCYm+m+WxUZtzTdrEGAM7LPvJbeivVOq8sd0wQmi3jD
O6DbrE7oYAFQ8xIHGZCFiAWo6h4XIsF18DvrwNOzsLzTy77D6yAgMJaYRHYv1RHvppsmQ8bkOSP3
ibpV5KTJ23zAzByTOTMK/6u1QU6scaxrJ1lK68TZ30D0bd0H+HocjfpwkaFk9lSlCaF5PkkjQRug
UvEpCzOjgmDHea339Ey7GQfnI6trPW7ReybhFEnFNoatSYQ/mCgm+ZWmbV86ZBgdtyevrDDKhSK9
bO7F/8o1kzuBzzbhMSimEk/p4ahNOt37F6OoO2MfSvLx1HYVtojDaJMTz+Dtle5SEx3WT+75uwpK
3Xt/rcHB8RLPtxLR8ZbGZsWnHuKW5P/sjbt98/nZph/aTB5+KBqLB+tfehDd4VNK+97OiW1XyZF/
Bkz9JS6avD838cxT01MbiUX6CBVmNOsoUFbfIiosEvf85AOliGLKh3rdks6xWKjfkRSGAA0oPaNk
k9YJp94Zkp2j3ISE6YNkCHhgY34G0rkw845uOBw4sNCQjgbXvwBw1CXtLeas0SicEL12gsv1G0ZO
LJN2JVlchcIV5T3oTwVOAb/aRmW83QoGQJZnsDZ0BrtJmCkIbqmz7eM20giPBsKK+3mO1rY30p+b
jC9k/lU5fhyhUcQpBH8j0hsCdA35f1ECcrIi5Ul3vKBHXV6DuN852/2tfRMs2+Tii0GO3SrCtDUI
A/VpS9AbxA+yOkhQoZOTs41M7J8vq0Sd/2x49tobo03DPNhJILTp/+i3FeHt3HIF+gRvZb5Lyqfh
JqEuXEMYeGI4gUpiURKSG4/489iV+FZZYmlTjAWzmVcx8OE5B3ZZuDk0jjbWW+Owm/fJDu3CA34P
JlXlNM+yUeEL+g6CXBIsSyIEDCmZ5L74aQpPOqL4g31BXP01GolJ9IFPMhD7TcREUtS9zVruE3nc
cnIHyb7/XC7kgGV+ZekoSKbgUEbNSM4qaswBza61muDNhJ8SsWF/ufdzGfyHGhzUlfqnSeiEccVQ
HOZu/NRg0bMRVrGpR92tKSGpfydfVO7WmswT4q+TBeUq+Abrlx3HndqIhs8M7opMyKQOaPznXHDJ
Q17JrpHA77g8bZafxuC8cP+/SGPfkVRcQTUwhsk22VYu88nFkdwneG6H5YkA8okeKKV6AxDJSIle
BkUtwUainWilaqcILQGo3hWA+qhIcyTVB1joXv2y52wbqVN5w3EvwACg+8btAGcpa3HrWZNOPiIO
/vXtAGOVc3KxUO1L8S3OudeUwIo8uckzf6BNjSVcivyEYMv2V9bt8V33YqzQva7qLKv/f2HPUDwF
QNaFp85cdqhQBgWNgY3QeurKA5/CAMKyeH4gUkuHLtElLSlkmGSRx6PwUMXgaAkFGYc5kqDZAwmE
66+9PRk24Zurd5ZJoAf13I8E9WE+6lkYzcoL4vnmq9qfSf3MfuVMvl6z/SkCF7u9nMzjEIiqdusE
uDMP7Yz0GGVfvYFopPLscgnf3vDlFpe0hKFO68bemhI9tDWFR+8Lq0iFJlbmeg7tN26qaOKBLEJI
bf2qdPA++L4PXXD6csrVpdS9/iwrveF1u+W8rkjWZwZqMhz/1SDha4uP9RZjUAi9Ahi54CXYMdZH
5qJq4TtxSH3gSBXKtQYXEQ/fKb1W2PvpgIsAHK326sVyafm91002NoFOuj7aEII/JkwHJOFyo/0F
7Xa67O+wSyZXG+IIeqRBgbddjz4l5epKEN9C6iFrgo4xhWjbzCnbOKTAkncICGyk8P1jU2/iY59h
ZgNHjSSS5+hUiVNrh47P0StZhQqmpURn2svMJP5o/HhyvOtu2bTQ3F5puo41ABk/l9/+EtK3ad3D
vp4F5fJsgh3KRITXOzzCHNDmo4fTumtrUCwEIJFifbgiQkW6+fb/e0KXPQLrnGiiY/z50D/4PKiK
e+nBJY3dAcmo85NQ+ktx5NUIK6l+mDtYhffnl25rkMjHWyFJYvT222HMm57RgCEqyVNuRcb1Pr07
jj16/C5d8bdWlRbpIHMcSEb2EkKsWbQIrZUu2mRrJIfSBYFmjlkvuotfWrWDJOE3wAdvEtoqtxqb
HgmPlSMDQoBM+JWJ6lPRgejA2lrjXjl+t42gBknQ3lVcNlv399fBltBUSOL6KY3orsU1hKgASaLy
GMp2ySlVObdlsOzbFULXeToQU0WopSsAqEMniamcebJspUlFatUKNAAwvjgJfHLkNiPKE1gPGMw0
mVoR6k6g1BXpVwQwut1shOTIaGLsHKfbDZeecHnffgleCP2xwP5VN1NZI/pDXNXDPMPXG6ziZ7KD
1GFy3/gnQA6DJPAIQod3xHQKpBfJ0amPYmihT8qJOvNXv/ACq/iQt45k1dWpGo+QYmOtbHM9RC6O
UFJcAQhqUGUJUW2vCv5jGhcOts12ERxcAUlnoiOwkZxAcEArMpEfi2ooL00fXMkWq6qYo9EXaPxl
1PJoEiO85fEXoEUz1d8/9Fpx47LL65zYAhx6l+DqA1DhxY2oPIBm4E7Ev52kfRtEDFfnYZNjXVTQ
y7wDaL+bx4WPnsxqvX/GyShGxAYhu6zJKGa+DdpfdwewcJ/eT7Ff09VgqzCdJWzEXnxn8Sy7ow3e
pVNl3Iqj9NI8nd6b1Q+vKLb1xmJmvgEYUnaZ51ulFM6HkJDPjmNFcuWw+1SJcHwKYttceJmYix4g
1/kTQ+VPmKyTKqbYUFFpIY6f0CCuUTdpIEUbtpTERtC1MgglOJKyc8VKSsMnm7j72MwL4xbc/zqL
XQtlS32JL6/kv/frJ/JngTe0+8tPaTKhpqH82AvRU4DSOEMkn4TmTCE9g4nsqqM3GJQ9hsYv03jL
18GgFux2Koq6dYpIOmWIjDbIS+sStdy8bTttfRo2Ye9t77i3v5sj33M7UXPxFApf11NIwvuUOMWu
OEq+1hVA8dbW9yMBsrfQGQt1MIN2F2m0yyMx+o6/+P0XHjD16gdT3ockbZHLfw19Yqj4y4BAcElT
nR5aE2r5ZT4kNxz3xz/kkBU2YZHgoYhfJmBydauZGLkmd8WtjsbGAHaZ1rwe3vgkP7NxOKSrNXLG
1giWTRDnqfxygBIlQ2LcSuKT5wl0cehJWuPJxJUpwQkHvm3p9JBJTUeM7R0AR/imgFF68GJ5lH3a
SEIsmFeEJ3vE66odtQXDdN9auxuHNJ+x6cNYL9DpK7HU8K4LWXgt77MSAcKMzoCd14Ff0BX0PYmd
Aw0BPEBQ6HVks+c+MSJFTV6iPnNXDvp5kX82e9m5g4hEKRdzhsEm+Tv6x3SIS/uUFqJUkDYm3Kz8
5JZ4KO3W9p6bDBeH26jZa0DrCmGPTzvSfPghLuUoElhRxGdPQuBFWNybnQxWxWNS49eg9KNp9Pem
Sb/D5C+5to4gbRTCVyeSBMvZQt01us42Ob2SW4VUz1psFaHQeSOBxV7mjHlnlb/h2KWWuL1eeGtQ
8jnJEZStBacpyNVxaMNPukmRkRlVaVfOYstwLwj1IDagmFEFrO5Qjf1Yp7w1rVsrCC+KE6w+wCRy
mtb2SDM+WDU0AYkCpuNpVigCoiuOAPSupe1YNoasLOjqoIoF8DmrTKCKt5n0A0VpU4/sfWz8wCO+
qyXUZD1KgkgWG2tk5mPf3KOmxikbOVCkqOXp9dx1cSA8dkKFtDCNV+Lj+St/E6T2htONJtayFRD0
waiugwhEHiL4VW30YV9kMm9I/gtQ42bVguCKCJ1R+V9wNqtlj9dM0qeqnelahpapq8W7Vz9u11mk
FDDRHQbfXyMxmlVNVNJshI77U6Rt6yysAB4UPGzPEZdUEvcWX9DHj6N0SPqRT3fm0ojh7ceE8ptB
XL5w+CaZl8BP+kIC7tKE8oxjy8zdMiudB2f3n6hzgrrkImGnaeE7W2WEtu+b4CsCby/FXND/DqA+
MttMM+HQKz91tUmiwHCYKBh6RMwhJfLje0ZDpwLVLnT2KdCKYWRamZ0nuzUxUVPf7q1G+qZ6XxxW
mKTvIrhPR07suwOhZh1jqQIAAnEaY1i/cfCdCKON8ObuqqvSSf7Ksqy/SSSPYFDClyzraaWMMMiD
/9PEqagupGJMQF21Oa+PnLUl83/rTss3fjIQfUZdCykWWk6YVCNJ/3PBFRH3yfrOZSZrsKMTNtWe
ZAIscA22ofq0W08AZi5QRZSGg1LYrS9FZC3nVsk0ptNpC3RzrXgmb47tVoSHSo28nH0vSznNWfg4
jpvp1qs4IxuBekDehzaP616kg8SGTJW7agcSJtbA4RC1ow1g38Gf5hHBQo0VnpGpHQPxZA9XBW2W
aopL1+4njJ3xheRBbqsREnv6e30pdoNpUVTopIHPjnUtzw0an35bj8yVa+eDtJZWOF7h1Pzhz3bE
noddl8kERfgLmJGngF0zzrVButb8tGKabRuvf+1lA0fyRqtnnbwvBZY//0pTOqRTDtTbWPSJoxvG
q61xfQgbmQeNeV8GwRQN0PfJ9tjJCKfJy4v34Uy908R9MV/poRJdbmYiR+wYl2NGzqotk1uVQABY
05kZNb5Q0UkrTrmpF4VOujTKDXE/8hs0JowM4OUUoKgmMbcFXHuuEwZqxdWqnOTvzQdCvYZj5JbN
kwkoKBSevpsNSa6ti61ax41EvETd1wK5+5v0In1E7dAL+832Nl4fT+O1+LUz+cvZHD1yLw5ez7fw
bEmj9lrfl26cFgSUWV3+ePcFrWvaz7DGofMJnLwrhc3G2TZI2NAnsFsrYnOBBNwh6avmBj/Gk5jc
z8yIb+ZMStZaU//Wt3NBv+s187ikSf5cJDBMziv2OObYATzBhD4tXRT96XCsCKTXgvA/mVfJkHVP
NN5Jc/SezeeYepNgHbhLTCtRKeVUXV4PxnTWPmrql2LtLkX35S1ikups8ehPr81M6c2nZsu7iwCM
N8aaX3SvV1tlDiiB+TzyeTm2nySKW6YNLuLTK37XWpNENjMfGroV7aizJuvyNfdoalaOEdxktHP4
cMCoitQpe71AxSRbBftfsKtPNBsmsyRmz/HBlfuuNkforlcWadEdrc+yMUPkMtLD+OqVL8uK6l6E
3colCrcRi7PyDAc2pV5mtCTXGQ8LgqObp0bHnGV+rFZ1VmP+8w7IloYdMr5YtbhfBklsneio31Au
JPusbmlCSJcWKXZ6BHjp4bS9w82/qYYtQWLnu6zBHOxpONiL9ZAZ2YRBRQ44EnHUMCE0qJ8SyQDF
z9rdOLLJ8NVA0xFvC6zylnUExlH0BpJK9ByR3uvMQg4451KOS4dfrD8rbNQwpH+MmnBRyiJxrC+G
nYOXJDHkFKeIzJnNS3f2qwHBAYvtF5KCWC+lutJIQEsovwhJSdff72POu64ko+yS5Y2Oz5fbUzQD
Z0xWEHvFtC3517IRudwW3jN+cV/mzSukYquJ+1xlszpXvl7GSyW60QHPdyBLxAUSklzuDnJXHNfQ
GkHFsUWP3DxtUoi9Q2KHSDigipEb7uAL1YYwvB1zTEif1MZn+JTM9KYcQSv/i9D04JKYPpRJ2Wbw
j4736paoFhFlZc8uSBqaXaKZAA22w9RajkaQkfW/imDHMmaZiLcEtHUx9Y+d7U6G5uXwkaTuDT6k
9XJ2rHh31y2aoXT9caALZr/Zl3EL8jI6Wk91DwjhKrdv8npUVoWI5iA0XlRjpa4k+znOUKQLfx2C
5vyBcGN8qetdVuDBuSifP7RNEuLYAtk0hCEUT5VGt0lg/hjlejqpDDmWcPA874aF8SWd+6d/NaT5
h1xGlRnztgMV2K9dN/zR2z9bwi6imcSQLG/CYdTaKZnaEUAOci6G/wJYmRhAi8ZgEkxw4/U9o8eE
Yqtbry+wX9hjiXqJM7wro+ZDVLYtp/XHOz/fN28TFHju3K6EUUM1KioJzlyph/9AQ2F5j2s6lW69
cCl7GUYqy8k6ROTwcJ+jpwhHOtVkup2SPvWCln6sVIgRLWb3iZjW+334aW4itGdA6Ot/oBMSlhn6
3nKT1JapI86Ky0tj6qvVuBeWO8+StZXCpDi5xixnxoDBtFiwDCujrJVh9ABzk6EIwblNmS004ojc
7JLT8/+70KZK86+ocFq92e6+cymqm6HRCL+B06IFpRBtk5K8sgs9e/Qr40jTJSd6zLMr9wp5zFsL
Z4WVRWKU0UkPfV2dK+3N948Y7G4FHJJj7Q0J0pUWDUgI0sFnAsjT47m6+oEr/Y1LDdDA/A2CSv6D
O7HC40bS2JptLZYZWkNKVHC4TMiSJZ8behefTgTD69XhDWKv25ewJ5K4EV40KLohxVka5eYHS+bw
PDtdz0ftDNDEnBfPRKiYjs+DoNjmED6ZZw0lCPhMpkWazW7GEhPzQT60Mp7g+uVw2Kcpk+fv9sdD
LqIaooog0Faw+e4Pxp79TZf9PD7QpMB9SxXRdHH0eCpum1b6Bg16rSfxzMU3Ijz7cNBrIj4+z5ew
soq8E6a9LxJ8Mk/NLf/jqNjqnp5d3UCg2qjKAf7589LMoYdy5Rq7Byxwaf14DRKEndxW7JadyjGR
mNl49DSFppdRshiWX0earSAOZwTYxnE22epo5U9tTU9NCohAhSRHLWasIecisr3U44YW3sWM5KZT
SmVjo1ZI4tHOahniuSrUZxACatuHgihpqgpzNTXu4gDS9gsxPC6uI/bPkQc/0npvGYALrtLB6WDH
B1myuPrK03j5uHL2R3AuE8/FBvx7APo38aZduQe7t2iRs4ElBh3HOLacE5TbsxchnhTh+lMKRmHH
WLmlLoc5mJQ+7MW03+sTNp/GScDkFtTAfOzXqj/bp+s8jHFiAndnTejIB5uY5XFfJYIVMdOxkSkX
rSKtteR+UK5AdYH1qktol1QD2FArlccAveBWs0tj+f3qjeXMShx+hIR1sReiR0c1BUCwo/egejB+
xTWplFQZ8jbE3S5f+W6G1z8WeXT8WvrKdCMAYioEYSOnkbOOtIuIy5MdKRTc5czZ0yUdVuCaB2Nj
jRrboypfncKWSVKPnTLmytmp1YVhm/Pupn6di+tZtdXNquWt/beHnR/LMzoC4QQvMM/iRxDDz0pS
4cRz05sN5HysP8KZCk4YJ7CLDZs5jldyyLOE39jhEP1dnGocjAnw/jYOFeCv8ynYDazq8G9kQ6Ew
UyF+YsJeK+b4Oe623ABY4iO6uo8e8QD2re/IJSf5JJaR+erTfffIoXlsR6V9lhdKJp/gyDegLFhf
iKoTQn5HECmxntMlb0iDjsxWTDM2T8XbIhBMPAF9y5MZ/+hnCw1Ev9FjgSp8JdVTDHVUhxf+67kS
TU8RZy4iAbJB5ygptcr6EhWgkZAmPAy4+NTOmlLvm8jMrLNaqFlnZjpykMf7BguqsmzWcvw5yR+v
VEk/6P0n7I8uzxB7Rit/e7gspG3a2s3AA1Y3et9HXg5fMX/n9M1VrwoKAs+z/t05rsFii+n/qcPf
dXcpmc+h1GfDQeHS8Ulc2eEpX7+gQxvET7jWMZpoNDBmqx3ybuoY0HaAaqf5ndVk97GCu0FSb+s6
wGs7XJrczW063izf/ptu4t2oKZB8zijC8+sDg4uOqXzcIS1MLoAICoyiWCUa/9A/dbrYr/eCUPdg
N9z6R6XfWALDWrdrpzCORD73dTWQeIFdnSQTK0MVM10EdkkZbFcaNvuvMCeGI+Alo0nKFskqKjdc
oSHMbR/ZeSL2BAjV1M3Uv0IDw9ca5aT5lJt8lE15LSURhwPLx+CFkinoQ9XHwkGEYjBS/DcWLrPc
YTE9In7jbLneH4ljlrBZ80iEeKTBs/8acRlCkfQM62EG3Z7r8zIjnDSBBqQz9itmGlNjT6YgXXcU
bd8U/ZgUNQ4Yv/BYg5PKmwkfe1Rb2aQ/AIl7WC0Mek/XrA3mhttfaWUT3yfJJ/ngE9PoLxaTAnPP
MUnAxJ+tY5NXIjU8Yx2qtKZ/HPrUtImhvVN/ojGvEaB+wa4Nd+klbAdCcouMs9G+VE08RN8XHHIt
y5OfZhIjoutBe2YumIeAF3hJ0ImV/zUDUqKrLJU8B7byuNJeoq01j7+dneixASmgygWZ3RDUcK73
PdTa0QBiW43PDsyxdkAk3mgykLoK763UJd8QD0jP4rQFTBFtWmQ2N/vaPQFXRH7Ecty0X0ZVRnZz
HggGBn606rc/PY8RFQZaAsnLM6KqebxHrZpRkiKJyveqS8ECLxJJoptElVphDz/v6a7IH4y9iRV4
b74tlHJdtAm2x7mVGrJ6A8XpEpRe2IcDtesRY2LJ1Sp1cHGauGkqBKKeCbjbkBDbLr10Gi1ssZ1P
TuEwMfW/C/dtHDuZxyOtRJ5/SFxwMw3l3+FLhsIar4fCl2ASd8/Zo3tR5ktQdBuN97RmKx1afMYy
QvxHZ3d+PDIajx48SJ9LWII4c6u/WfzUkA7AzKUoELbq7z75rHXSNI2tymKO80GSsDbN2zw257Ch
BQoRWmjX0Q5BacL5BvnC3PnAgZpR87ASZDAsQ42awl/KK+lzzCQxDVxjQWCr/b9mnPBjNaO8z7Kg
S0EaBhk9BY8WoibFI4lQ1bzNIqHpBQgchGMQ2fQ33BKtV+nIhHJGwj27q2nP4bh+HzVLyG8/4RDN
k7le9hhVuWMrtPv0KEu7353/qoWHdXUIPpzjGvovZACSaevBNrt+DtE/lXQDGiWOXP4hmptcACa/
S1HIqbTjOvCWx/gw7K9sYjWDX6GPcELWqBvtIzcVpI8iUDwq8p+5vSnvjMvNFUkkbgHOLfgDBO6t
Y4tazaY/dj0akemJ8VKjjRmrFKZ9vbA1z6Cw8C3raf0DnHBHWrGIMayvwyI5DV4yuJbZuJgfNs8D
gk6XGDc3czxw/ik2mTC9lN0nbsB1QQR2HStuhqEKUc+Csvh2/nDkd87U3VyiBgX3TFqkeN12Uf16
muQeald0Z9/9Ecfv3QKntgxRhXsjC7kvZ+7vqeIEffBSDZPEhyPtALQlVDFfwLEbvg5R9sq09c+H
IKXb0JHYbkBlnrKbPsrblksEhPQq+JdyPu2NdDmkIUILwrRJal0GG851mZ5OWAqsOKNlNcvSjpxW
VfmbKfUQf86wOI1m/FIhRiI/Q0jGnjc9i1C72oojXGUA6OmR1om88HoNkz0t+aGv9an/O/RNAp0A
MHnCLwLCLBCNIzGfwqzbVLkDMSdIeYh40SjXUMpZE1ucEiFP1rebD+gjwVTlG+I0xa9S1WYtwd8C
IPsr19+SHy2UluzDuxN1oABPV211hONdq0/c6/IBCJo6MSGG0coIAf6Q2R4l6hywMt3JNYdrjWEU
iT5wymyscruJItPZbA1px151r7nPXGZh9VU1sUnFfW4psCY0n+ENPf/T5lcNQ+nx+X0YEMsRGsMg
TOtL0MAJkuftLjnELzUv11CPvwAsV6avO/YX6KhRrIoLQSNqoXrlC5DQkcWXQXImDlpqaS3NrSbS
9V1HsgzTkh47Lf/DDZ6Z+akAy3O9xnZFJeeeIY61GEopRPsznrr3RN5KO1R9lrzBPudPGbF06Tz+
vqD7jSJBmCsoHYjtFNguve7vR2OaxtgSPrA0mEbWLz3oYb4h2INw6+6DXuN5gVpOtQVnl/5Y46RJ
QLouebus+0a8ciUPLxq8XHylEPo2U/C9Phm4v1bGAfgoaqWBejHBeaP+kg250kyj2B/EA0O/gcX8
SUoV7mdv7GrX558tG5dVVcG6FuZLy5uk1tIqoEyeiejTVmHgIRlEI42ItdWMDj9ay+uXZE1rJlgb
gA48SG5F8mjNpuXbbJS3cKA/6IzmQ5JJxBXli99hWPuZhWWZ2mfcbK7mae2AiAib4NcrtMjRQ8aQ
zAdCG0yMkpA3vi05EZSxe+84pk3ZsI5t1+vI+1Fv5LdzJ8zuL5+Qgae0Z4wDlOR/Z8OY/uqsk9io
MdKa9nPOmIvb+y4gz06wRrjMd5+U15ipeKdKQ2fqR9+wqXzyXYzpipeVGwOZkxTFomJnCzIBXADm
YCl6vIAIDfzox6yhM5lapcJpG7wY6HbwM18viJ88o7pBC9xG72EQtPvjiK8100jkcL4Mtz3lFg2h
wLETF1/M0LzC6Sk2CDMbP9iqqr7TVfZLuRdIDRh+c0l76dak8ivhpWSBauuRNUXOgFAha9xV8dRP
21Yxbpd2ZCjEV4Vz8LA1xTvi6MQyKHpedU49mZ+JQ89fvJr/byDR9rwq0XcYroLQQz+QUkExTxe+
hloDXVqS9VFUJHxiRKln8IcERdMOVmJ59Rwm+XO7E32qyf9LyktCatsCGS/xBhV6UpiOPMlJrNPX
EQaUuy1evWUVDdrGg6aEUCADT7MIZbUeFkQCEPZEFvEO7xzW6HRy5EIlZoOGYcK6UTkejUhFGvz8
6jOh/It+E5o51Jy/IcLCTED8gMi33g6v3qy3t4B+9P6knDTa72CGl24c7S69Rzxm/F0MP9o80j48
zNuFwYpyII/ZxLTQdPbQLzuAwOnEXi54twWdfRwasCQ1N3wxISxUkxR/ci3EYoTC2tZ4Ry41v+Zb
+s/XAQ+qpU71YCK78ZJerlI4f0hdAkbEDK1+WSS+CxASQm9/Zdz2U2XV8XU1/67XeU57KZefw60R
RiY3tBJOVhV1+4nsG8t1X6xjs5ufnitbKha58vxytDL8j/1oqRqmAvIZai0jcksc19w5/6u9ZZLH
tWTtA40XyN2gPS+OsRwfmiyBcOi9FJK1eHqK7IPUW/+Ft7SOfJrJG7VKtoLrsZkVe/SxMNalIk97
faoGLICJg55C3Nkk+Z7USC2gROpvUWtqrsrYIxjn8Zj4riW9H5IC+1lgDOgUpJSOcml2RcAVC49E
6z5QxuCCWs5h3oD3Q5ILrwsqbR4RHkrWIPPSQeERNvqmI5UXDhMntWH1j/IRd0wu07VfceWpElHz
31WR8Qls0TKtlyK2c0gZ81TeRuQoVhwJXyUwo7JzDvD4Kx2bEMDyQhUQ58j6IXUf9cZVcLz7thJo
PXmCqocYqN3qFPeor2zgM+VMXDqNHW89/zLZtSgaWv4g18r05gCA4iJWEczQPheTqXJTtX806SXP
pU9XA64fxeoPBJZTnSaPOhX4mQFvOZpqvPP4Qwylppvfz3v9Jo1Z0MIuzB9Zbg+RT2aO5N+voJZv
oVY+NKSDIFJmsmSsqqwXXqYUOCHGCItW9ej3e09P/bhkAkqEVuMaIv3fjGaAn2hxGrNx5k1ryLa3
/Wdo61ED4ATXlaQcKXrYrFI1aRWhfxgHKU88l7pVO4rwpnheNSfypnabjD4AGKMiYPsnkilB0PVP
7Z2LrkQeF43VemUFpL7S5XmqCyXxkYxiHyxIyKB0yFi0EjPRGPdFo6ELWxAbOSbdC4jZgdqOqPVu
aX8ndYq8ZryfVBLVjt4YSXjr9cuIJpnoFI7le89kAWa6mwjXLNXsvr248yYNZI1wqnubkckj5DAK
0mK8X09/SD/oUYnvDYjWk5G+Djtlc7DNYckRBxUrbJmF4psu0szPcEWgBOAd06pARpJJ4sTL9Du6
nvcITHwozv5EwdoDubwbobQ7zOSSNwpyYVxPL0qISWf2VRQvO6lEhBzOK+bISiLDMaEf0zS8JGb1
hdylSxz+ae6J6z9NKX4pN4lFhlcK5aYR0Xg6eWRFsY/tyeiHSOwbXIqbSE1J1tQ02bhY7D1NU/S4
A1K7Xw3/woVKZBhudFycQ1gHvgH5EeXjRsEEYfi1Vna5HV33lk9w6YML8G9yMSzlsJ+YWYqe3CJn
dT+XSC40RddaNvL43B+/UVEdkZx4loOa/GICSKxa0sPOLZ3an0JpJezhG2VDJmiLQmjcR8FgkY19
R2BzeWLi18dd0bVCpuMPOJc89333bGXE01sFs0RN8OIXyuiWdQIg8MykzUMvKt8o0HNxOto+Zz//
w6q2P1qAyyRHW+67UO1aLU8d39BjxW15DXGJ+s+1RyyCJ9QWiF9m3udiJSTJXCxNqk0J+igi9F0R
dhdz7wHUgm7+6UFkvjfxDR4uRbdmaEshVLLDkJElka27LX/59dbxYY4vBgbC9f1vMXfxvzjS3a8U
1W6N13pgyTe+KWATepOj9SZUZnUarfIdXq0+glEr/vxQMqSpzoLWpdTYIiW3znFW7BOtJ2fdwNWB
OtQGJiWPQKNXJbIMcEg9zNNBZ9XlC5BGcVAoH6nhQamau8QfkR/6ZDa2uxAPNxgzVLjw3kxfgNL4
fTrB5PlsffseS6XXSyZGXV8S6Z29SM5YgFajylZvVQcHI+EkvXAE1huex2PZL29NTeMERqZlPQUO
gXrtp4l1LebGhwIcxfY95UeUHW91o52hSB91SwUlggSLa7ouftJ1LrPq+xGKM5koY0+ynw4/XAPs
SUM8zLq9teY8z7ow+oUNXWjueOY95KnjgrqltBUouFVr9esNaMOv8FdCGdq2jaedLcl7mPF/9luW
m0JbTw5BgdvDdwmJwxV5vCOeG8bPbvFtHYDlBeYuMYqrP/d53+YD9tbUmkQ6oWIVYTdPD3izYF+B
vDBcBg2ceuYSs0+/zkwgJlBLUqjBxtOai3J6tlmSg3pRrFZtUcBAlr35a1PkaNZuw2jEBUa6Eh0K
wtH5vOiNktANG73w0b5OiZL5w35Eb09m3GSV4Pbq95sK+8DbVLMsiYtQBiaefeFCHpND05IkcHRh
FWmFR3iVBwa1ekO1P9CNw/uAaR+DouTyHobDnCQrov5LfWC2Wk3c4pcS1ABqrrxmZ0PPvWLRo3Pp
h/FsTAF6sKEPw+wKP3rPblHi8pHib8O07+s6C0+FebE2BCNCoC4EqIUFx7Ymur6/Hc8NbAdfaj/j
iCSqrHffyZ6Gd9LNdkwWbi/9rbWKDqvUlgksWasIS0tmDOPHvN7xv2TVAdTrV884TIVW/hlTi7z6
wIJ8QSINu8zCrB2odWzqxVbuYpqXyLZMcQgeOtPUTsY5TndJys5fLR0av73OsCc/nexv7xwHsGM+
QwXVtq+NNDCn5M8bog+qliUU7+WY/sQ+gOMIv04d4ioMqiGtQ9NrKesRz3b7oIbhvssy6G0tamtv
oJguw9FW9WpYvTkskEr97VdpwE09VNE4XBZ2oZyAZd52ROnLYhTd4eSiziz55GswIfr3iNjHHKdj
z10j9HeY6B3aa77Kv+pUybSsA1D8P6zYxHgFxLgWUYnA8YJTQWRB5LqRPZ0tla488nP3lrSGeT0z
2T9B9q6Z9dNsUk7hCpE5/vAMuVLPY705abO0WawldaALsezY/D7dKahi2i0Dcr+shyNytyQ1Y89I
HbjdMcBLR5cM1uNOZlEL0GOxKdMqAKMikCOd1dXf1Blrv1sArKjsXhqvmsGfVhRvVD2+UdP9E9XQ
S77AuRd8Cjwi8NysXRHVN/Dna4zsPsYaYZ9p6TFS61xAHRRrdPz0+4guCnJZdc+tIJOR5L78RTzg
FaJ6Dy75gaVm8LX1cMiOWEdYQpYZba6uP6hF4h4WSErg0wLUBGqLj1q9WqFGzS48ZHuws5BH+EhR
Ul+cha8MyOXsu+6qc2wbzVC85rOuZyOeK/pS4PJP0pmmMEmoPZ0wVWJpWRHFAwcN8KimdCfHnXUm
8v4EyYS+YG8C9mw2gLKbZQjwr3MiA0ycecXWHa4msFFuxkcoB0kJPw4iWLTjW+1aapTTPxorwflx
KrvtiCGSKO9v5q3K/2sCLNihY/9iKho36pyj2ILDr16v4CTT9SHOV8P78ej2WEfEXyzILHoyOWNy
pfIZxgtmbQwz96QXz9fk5GBaJVPHR3BnXQTsxAshqhPoJgSvEcm86uRhk/lcfH4uOr8xCmjZ2SfO
JdgiPilSuAhzkEJFW980JqUJR5WiQJjBbLgvXHSZJxwmwRv+DEWoKcbumsttb0B7wxWd2iCTerQX
lBactewaj8xfmWBk5cOXp0efBDjQsLqldmAxk0t1TJv+vcitE9ZiXweaXFUEOiRnmLX267OlPsbI
HnD2faBUsJNoYKhReUDozq3cSLHkYsPtAUA7UaK6Ggt/GrbNYOWS4BuTmWGLL84EGbUx4mL7T6Ib
x0qjqwmc+Gccus+7qjeFxQesX3+FCBBnHZHaZlHCOP3Am6zzLlFS/QPHlPR5UR0TL6NemPy0rPEq
vupWIL92tI2myqOUu07CC9SS0dJY1NA8+yafwY0p9XzAm1CJQ+EStrgTgXzfNraGJafIXSkjPZVw
qBqD8bra0RBAOhiUuruXqZZB2r2p0EIeIza97oJ9pDJ1k45rlyyRZ4FWRjOiK42G91OOXqNkqkMp
CgXmiCfRi+OotDfOUuU3OpVrPh+0hAb3eLqtai0XG3LDchfjVIHtQwQeVZwfV87TXI4jjP7Zhp1Q
FQxOXPcL/AH1DSzEXfcQhTm07TYdzF0pwtnOXGX0r8BqFawP5TAntBah4jvak80rXdvmEETkelGk
NF7B4C9WQvHPVIVCxcTb3kMLMrpaDGCVXTrDL+lrIlxuxXQyTpQHgULBMePIi94Q2UNCleydIHaf
8lPFo0/6m0OGFBApCPQQYbg3jFcIIayaurUyk2DbmQdATZu6tCl3wdqq4TrdIXSLCXWfHpiVxYC0
fxepdt7v+2DakPKoDLQBeKhiJys7MNobq/Umfmk2TnZVXOit3ghWkDGISrDrbT3dAqOvze/oP6bb
uSczGKMIzY1Imzw/8OahU8bSlMoMQ5Lh+KfyA8fZBnKobdpJdTRyfXaUjeH5FrLhNa/7BHrHNmYQ
Nawj8n22bHXV6hOmwmD4ircGYY7/Xu49lF7EfjL8uGYCAICxKvOO5YtXk7/XFAvyDQhlvvdF+aGX
r6VrU/N4bcORsSz7XYa3RMLXgKY2m1secv5cqjKho+6achcVIKxohiLq+1P9bb3Vhz8SCPVotmRf
x0y8CmpIUH+cbsh7un6B08UzksFqAZJeFv+1CYKqL1kGWFJXgKrDp5YsDXYRBfLoeuPul5LmWe6/
xbPnNrLC5FAio0rUIxLoqNNXkrKfjDpDXWmyHJ2n8hyix9k53+3ePQThqN/K0dUP4OHhDxZvmd1M
k1Fm5bN+syXlulgIz+jYVgQ6mkFa9EHH7/fmVHsZKVNj6WCYtnuKM4b21wNb7DXW5Vk8wzX5fA7h
g9gRi3hXZ5+56dn+obnsCsFpuKfvpgOvRD00qKKVC5A/QmcMC5MVeuHGlRl3r4JV2BUECIRxfz8E
uI7+/eWczYVdYwsoinSZOnY+W/szK5C9hsBDNenH9QSnF9qqFCtDeBpBLajvVAXuRwfhDrNO82c4
IjqjiCVLN2Q+bt0Y5TyDGrOrsRylQCPRjlXEDYgDOezZZ0iqRSl9YfY2gzQSnT0p1eFWpcKRKG/e
EE3yoWC3AMnQe/CZZmJQzzxt+HyaDYodGywsQS0gL1SqwPKEkTLXwToos4W8iPi6JYmmkn4m0+6T
6Vc8MOMep5SeR09GMtIJfzJZ8E/aoHAURALBUxbwLZvRDILYmo8yoJEsHWw0d4rN/aWhxXrOnGJE
EIsLGjdcYPlcyLfTCuP5YZuon0V8hLKPI+vvBRkxOGpsUp1V5IsdSxbM9AlQ4ITu9TRtXFvlI34v
FU+WlWQi4hTy75OcOHVCSuKV5iqZ9FrbxZZUArBv6DBR5eR7BwIPPCj97FGmthV4YZg/S91ALJIp
lbjhr+GjC1qvVzJhL8CMll3F9cuNedoGTQtBJw6IxvggRW9SKqvaNDH1OkPsR3xXw/yE4qolEX0T
cGXc1Sxab+E9MOtBqR7YZMphwxKWcYqS2Z6h3incZSNmuwN8qHyAOfPzqLD+gjfq0eqMUlXaGrgR
P8vsn4MJeGwVyWUawM0mLLPpac/3u1XNPxHLfDQ9jTGpZPv5jmxfBQUfbkaqfm9+uLkqK3zuykJ9
5602727MkPZuR3tiZzhBJ1rNC1SrIZuk5TsNTIUvytQbkwIdlHNDsij3hNHh8JhImoKA7BJqh/3F
qijnSB6tuIeHYbgf/dVzi1lOdHD+aCQ1EQ7cOYASS19byj21e6uIO9VYym78FGdDnsJrlsicGVcd
C4P2FqK2e4X9J/Hw+Fni1033mrb5JzOuAnHszamAY3xNiiYi77VMvDyNDMlETrwDr9bMKIp6jXCf
AKjtODTaQLi+NdIvTW/sSgdVNY/w2m37rm105XQA+CcjkEnmxZf/QQi5nHyzCku6heC6vK52/Ard
aW8GsvXR8lImD+4goSSRMQPjq9bvk0k7dIpOGVZG7nMQ7nYotuqzvRLIlbPnzOxMpulEfL1K28wU
FOK9GWJt/mISuAQ8cfcd3bh46U7VXZNJaHpWqpkcYvQ8jfj0k4+v48CKAxLf+oa40dI0wZEGczSo
fElTBFgYcSmMKufSoRQu0oFxj5760L0Bi5MLQ4iKtDs4/SWa4+mDswd6tUWgORDp1qIl6eqMM6WN
RZa1GGARL12i0aPQXIJqZBxnhEBq5caQWtN3qRgRnPlvxXAAxn1C27CiW63YQRTAFjSia3EQqYGV
YfojdzOE0N7PQtAHS7UkkauOz6Bl0XI46aqZRETGNrKxIj218QWSpUCzMKNBIySC3v27ipGgWvn1
dlm53UgkpQzMO4P/sSIbEcH6QWDbpW93JW41l8YG3/ZFnf3GQaTMfpKLCi6b0L6YFoPtsxtai/Ji
6DtUSih909WR7OmIlZbnOcPovfiMdgpGBtZedvqOnDU5QFyM/Y3Eu/74SEJk/BWgdkPD/v9T1GBZ
OKDmoJR7zPWHbNED1YZZlq8h9hwFMX+jj6/Hi4fSPMmyeLp9zuPMk7UZrkrV1z8PYOrX7sMIx8BF
KBFHLiwAC09UEkU5pUzqho1+lWl+cFdUVknjPocZXFk/WOuhUmo+yLcF+QIdfB8/rqbJBkYOd940
CuE9Y0kGURqCVCBXOm+XXaol6qAU/fRg/RGX/0LH0vZSt1L+T1SnTs7ki+BxAEI10C4POz4JhiKJ
trNGIXayaOtyxL/s/wrwc1jJR0wYcvUezhLQuyRGfS0DEbeVXpoOS0aHiMJGq9gdQkL5czoC1AUE
Sq4AIhwVxTWuS4j2gdPw0JUk5XpGJ2jas8LDoW4peKS5VLcICWXkbvxhjQU1qNZt6XEuFRDNqHxa
hdrPLCqiogaF6Kpr2HbU0k4Q2M2UgHbZmj0/oWbHfNKaojGMluqguF64FGOKCWPvM5SqkaWZOfw1
ORr9XSh+KTbUbExLSGBa39QHBdaoNBWxa8I/lmFeY2fGNOXnKiFzLmjXMiurpDaIy4jlbh69ZJlf
krTbebf08Yw28G9BAsZGGRV5UfpIQSLb4vh0KZwuL/mJ2xdmix66lmUDiG52oRaSHsgMzc5IUuXQ
pdLC5lIPujZ7QoL+TU7xTiED4+NgPnvWZeAt8Btq783vdFu7DPeaokmjhurqjugmT/HaJ/m2TLwt
0/hthYYG2zKEB87a6Yv8WE6A6JktS40wsw27Djgzerne2qqCT4uyt2wRTp6P8JdfgoLgQ1YgEoaJ
Jwbf+cYUnEn2jIJfYVU4nz9nILMMVaEuCIbnEulvI/6Zvew7s6p4rDBMHAa0APBNNQAPwcvr9c0K
LwzQd7qwDYKJW57hG0MNduQBoO2B4sPgX5FH2vnpQTMirId7wj0aPpRR9sbfLI0VcQ7V3g9tX/q6
CAk/6uzmZhM411G3vXbgoaP4Ll3hVkYz/cb2AudJhe2pd3jwCp6FU4ojz8T0k+h3QiIfLp+KYweF
cImzABY+4h5zHTXBq65kKaSn1gBMz2QfWJ+9tagbYGNtUwMVLFaGTJmer4d3Os8CELUdACVsKcu6
zP+z0ZCn7leSKZOdbfoYbTzjQpdP38bcLdj+DoZXDOQH/APhJtPgOM7VQlGHRtv97/Yr5vahMMlG
g/DQzlhtIRY9JCQjwKPVw8//aJ8G3WaPzWW6lM7BlyeUdZpDmj5c6PoM97TItMCjzTEulHZTPJJH
9Pcq9mjCOCiwHoMErp1AehX73h/5ZhnS2UBTDFqBYhfX3K46Si2ekzK/P1uAjwt/20TG5xuavuqw
xh3lV0pTIt3WDH7Wv37K2M3q7s6F1AC1KJCI+i8u9Gsi52q8r4Bv1cpgiSKMGJsxUUPWDgb9fF68
2f6FrSZuLSqpcWxg77zFuu93gDIkHoxAk+91tcuZHCE5apuJVec2VU4oUrqDFw1LVcGyGrhRJQha
1OtxA1qtu91k7Axj/ILRUJ20E+eU/TUJHfP1+BVYCCFnLcoc+ktX9CPDXnw3K6aoPRsz6xzbXjMc
sVCWtePrCZ4+DFmvzHLqR/KN77xGQoIUKnPhBQWzoI8icrRqmlN1NuLKi/9YWnF9nEyaPig0RJXm
n4cdQwVLNy8CNyzD0oIwnM2PY3cAlhM4HTLUJ76prW/nT5q58HtnyUQayNEYb/KPXGLxLfUHuJG7
9XxAt7J9fxCYtJYW1ksHIGCmqHBVK72jLs4eHrZzVEYCusnd5mMdTCJJ0XDZtp62nAuJAQDjOwRw
SSaZv6sAMZGfvBk1SeIM9wGIDNpNZKoZWZS2KwuA9DE6G67Kb6o/ckb7rU1O1G7igLsBVBG7ZSxi
WwnSnctDbzVJdBWogCgiiFIr6N79s0chgcdvo+kR9eGMFPOin0+AsvECCm1ux/ASHH7TI5er77V5
KoqHbNimva5xxvjZwo/xPwelG98MRj+d18A4BUKZQ/x1ULVlDAu5OWEy+ksjYsTDGU4A6Sg1xcRL
A8a+CX9ztIwVUrtNLtRShEWqv+oadM2emJInH2s+0jORRLaCd7i118wo1Z+HhY17CKXIVAOFcxz8
BMVl0zXIF54GN8I0wPI6FsiZMJR9tf0IEzBAbz01JlH+KWFeWOW9ROctq15jHmRe50OXlBWB+Yrp
RsV+HC125jzdCuzBejdMOR2YoN9Wjcdqmfd32hnpV1GEa7bsRhBqPwVa3newxfGsFtx3hynSpo/4
3OXXo8DW5K5ONuqsFI3RYonndHQn6EvufMN2jo1chkgNuR28yzuoYu2ncfGfAMgzGv71YFc1i4+T
OrLUW86nsRCkDiikTa1Ph9h5yzdpe7CDtQjuFO6AvJVUr+KesZsKcCHuqASfQcNvt/uGt/Yb1O7u
SEZECbmmpmi4sKLMICosEkO5niVZGYxGmu2bY76fn0DunXdVuWeKPFNl5ABDfQN9U6JO2RpFKoKf
Tkn7g3PK1wDUtKd69PMD0cHOU8NEo7p6EnBRVeTlCO/fmOwdmmly05+KGeJpASWur9b9WE+sNPui
mB/7Q5a+VhBulxECVQCSW6n1yY1aEgkjYQEJo3lH8jY56x586tMhtNOhNlvgHsLzsYoCA2DD1p3r
FiMwoYOpOW3WQ6uRPqBUb5SwgOJPPmv/PRMWMz5idnl08xsLkCdGqiFbFE3OcIkDC8Xw/yqa+2gW
eiAKHRtMAcdx1lZ8adxTviqBM6T1dZqJxWSlecQM/hvBnrhEXP2YyLA6SjxLd1HShxfqfPPl+6NI
/JO6RspZ7/JXrGsmaAWXKhaohLYhPJ4wuIl7psfcI5wkTzPY57zfuB7qZvDJV07gCdyJdB/mu3Xh
wknXYXE042vqPcKFeFztJ7rCiWw02oV2hvGlYoUiHvHtZbDl5SI0RhysM1o5kRXWS2bgvwzdmMiR
K/b6ftEAec5m2gTctWZiBsfo6UFaPV6lTRgJYf6gxBvhdXdzsqh40N8cSCIm+t+SH31iRyj+dlTW
4JjPo7uO2uSeyMqTK06m4fc384m9NvZ8d48s9yj6ZE8UynY7Q2aBMHqeauy+iqyYse1I/+AMmLcl
qaYQ3diWmL+DyODXI6BzgRP8Mts9Wmknb5T4R1HQwFpWMOEU8kacTDY14D4XuNHRiSitISd/sXft
BbkDiCpldgnr/TsJgJ7cyp/MKGhZo7U0bhHpm4+7h/EB2DeGVDY67X+wjdFGkvy2svOjmNf1KR0c
R6eILZkJxovKsNZcRqdx1+v/O6ZFGC25dcpyh4OCOQbBy9dJqpEbhmgsVfp/frk/JhCdMnHdtulK
dfxedx6JOU7lAKq7kspRhK06wgtgIbx4en+glqR8NRj9UtROciAyf2dYXmivUJEnRbcnu6I0eE5U
JSWW6x2Z2QZ5AGI/N/PFZngu/3jYFyzuj9fTnsiQZYmuE8IF7oK9FMX6zfk8AgBYg+2jO5BPO/PM
R57DwqvY1iRoOSyiWpSqxpaIvF06tJAEIAZ7OBru3LMICi/DOAroAEIKEek4hN02lyrxmxX+KJf6
WIkhr+gVzY4V+MeXO1QvUUT0ZvG6G8+maoKe8vVJTU7rT5D8jf9oJ3Nd+NYEL9zl+n9jS6/m0NU/
qZSmTJzvb9+pPwc5/W8D4cCaXyE/iwDTuiF5Rx8ehFoDFHQi+NAAGbzCE+zPBqKTLvF2zfcrLb2M
3qv8jNi8Xdmm2+CcMl4YY24lj4kl0eeNfPTA5x9nSw07iiF1JyKdhRn3Bi/L4SEfOTiBsc6RCsVp
45jUEfcpC35riU7bEEziRlhuQqcWepAtUvBgIkCPWWICTpMvk531Lf9tNsygg5jWCoPpK/VeacGs
SvV00fdnbrChVvzr7q/7nVGyt+zp4VqMpsmn51oyfjj+vnyH8YbGmOJauwj6ySjHpy0P/oEWQ/J2
iPLtP48JaAq7wYkPjXXAC04UTrhB5zfI3HeBwG/kO8Y/YDTZx7SCaSrtuW+/6YnAMd5wvxIMxGss
1KCuSdYK2gzO9tK9venZ368U1g0S98fSBCc04Rn0m1zPmZLo1aNYJ1weZRInR5DXMwyp9RbhI1iu
20Ez2zwscAnzDb9PaX4P4oQF80fvgnYOEaJjYYtnEOWYvXmc/5UcVdbi0PIS5xJnk6LCxadR2PE4
4dcAO6QYWXtPYiQIfJgtGO34YnWfGCUQWTKy7hH/+lK6GNXCzTyiS2LbmX7+wE9xfj4xvCJ/NIWa
cQnX93MJxhBOK29zdtBNHr7x6R6llqZMVsR03bd5aEuhZhiPy723G3HVNF07A/jLC8WKGvxx/mZ5
X0MFiQrGDzwWYH+0Gj12Pvc8Ud/vxFBAeb3XZG4HddYQLMjrHlXBmHTGmdmeBdf8jbLBSWl/vxw8
pj05uIiMOFXT7tPU5Gw4mu5V1t9958RN6g2H2t8eX0hgr+wfN61smfzkvgFpj+6NLWV5EgR5hHqz
iTYteVhf17A98QdLvSacKq2w/HQZA7ciD9LF37VASLHFDAlNkgcP0J8bFUeocgg9u6faaKXvBIRm
b5J4u0irXSG7NW9WzjV51VIDaw8JPr/TgYuCKuSj3MkU9+4wRvHb5LXLoWeAwcX+5qktGVXwcfQ4
SQcRBa09xDIFkLqDRL+tNiZmxZKzFQeex4IAlOjPeSUUj5BO2mrt5TL0GQ5chVlSTZMIgJqooQbX
PcvVSKCVhr0OV6Y6hCM3+KUwVkE4THI9EEYjf3C5IhC319mpcmDSQT0l1dnHIUrRrtU5mCCqe03z
FUUw68IbxSRMo73Cc8C34c2eEn4OQVRv4WrIeeVprkH/B7CA201nOoh5CW0ABIMFIuw/4Io/ZOyl
sCaxUBdRMLCSVFntPKkhUFtEcBkYq5vpXdS3tdrqv+zg23gRuVzcJqEgRt2HXdy6Rj3pNHy7AALv
GUs9eTNGNfwiGoGTWwz2PEFPqEZwTyD70xVKJuElfuA27L1FThiibW1qrFKwxTn4R6868HKFopBt
XAReiMyFvwnAjwMIuIsrlWBDmzI7tgNk9cb0H/AegaqH826uZsVBP43UAD8Mc0uiLEGEJBxmevVj
JxRkv9+k7qdgSvVtC3i34uO1avlAzJGlYtaCixhrTBvem2PX14EIwCNXDjGfXg6EgqqSqsxRfWpU
FmQF3AxivCgySBW7h8+DcnL2iNHu2DPVOZSDD+bm+KpQPnpKFDybES56AN1LyguXW7+D9gXp3xLB
CIb1/qtaUTRYyWGb6WpFI4jKaoLI4YGl8rVxs4lUiUDXY47N432g8fB7dje7nWCQ9iTFsjEIYuBt
5W7V+cRIEvyRpCL4ukynpajheY1Auh/jNgS1nvrudMq+AvHEWRAwX4LY/i1ggV0hQNZbnk3TeBkA
gYJc27sCksuLD/RqNlWw2NOSoO7xKw6iP9X9UeeU48A2FpDlJI+O/eZbLpbl7pHBqNczHIwt4usv
mrGzTGo5l5lZ5PNk9NeTXSLZTwx9D/gTTdfKwHN18m00DmN2krDDj06HiPjHi8y/+wtMGPiFhmxj
/w22xx6kTCnY7sLtKN1RoSP3XV4SMxy87Lwn7/Atlt5nfoqvjTsNXjrDsafufRlhGKOL4U5DYfrE
/uQ2y1hYwlHoUsKyqOlEfH1dIqRi+UV6kRQ+URU1wOc6zLan3BkXXjuPWCKTALtzeZJQbCJfJ+Gr
Ty+l45k7PNam6oc+Z90grjMSIAvCSZXOqD2OwQGPNOR2hwZH2yhvV9U1zdLG65GUPC2s38N2cH7H
2k9c3j9loKP/+dHOq+6hm6ojxTEVq4J3S5WSiO/gbzkWTkjh6jvLX2MXiT4GITE+xkjE/DGvRUBA
HIapTD5aUFdQsYND1IFXtGYdF9HjCAs09irUArIniGebB94g72v6rnfJEL8j+kbllbXEkpPbNLB+
C2H1VxqdhboZRHsS0EBKwMDldsInQ/shbQcE5o4YfKxiVsV1foKU21hfV2TByE7ALpzUtVEShfmy
VqbZPBYZEuh5l88s6IvCFk41IxAc12QUEnaQosJv5qrzPw6E0egmAHfZxJpJMigEsGCWv+A2HVm0
iO15cWKyym16hE1sjklYjBoCqZwtAn8abh7lqYttZWNxVzs/A5VNw/W5EBr56KLVPksnkFD3Ou7X
+TwRy+SKY2QxnfCglwctHFIDLD8pa/96B/Ml7qsWULW3GLf2lLC3Krz30ztufLCAkGklngBXMttv
EoAp5jhFpqVoo8LT+i/n4jE+8uIZ2qNRo2j/0fDQ3noaGmEAq9CYSTmC74WyoYODn+cVNYrmofTO
lE96kcmKXatFixPmI7bVyRo2CjLqIizK27s2E6tGpNof5W2/nzmeerIqHTj8Jb32G6iLaPlh/gk/
vVrt0Z/wIhz6Pm1rf+p7Jv04ItWynub8HMrrRLhjDizzu6rlEX8y1bRL9ge+HE/EzhZh/B12OJpX
4M5D60Ee43BLfbd7HPI1blFtGlc0r7e4QA+j/oxFt1hzNUfP/rigdlUOIt8XLt7nHl+U3aD++TeL
6OxV0rDwbPnmMIxGgaT1SpHK0KtXJQJJrxkLGSkicACUVnXEWJPAzgM72gfX4wF5xsdCPOdlcT6r
rdJAZbbwNd4uIzZ0EuDd5QcTqFABKeI2ELcvdOt15Qb1R51rrx19SBJjFocbG0TWjqAmtzN9Sptm
F2/T1atQHguFSKKPSaGJ1Si/63eLYBAtaF5dfBDVaVDHVkZHnDsUxmWtg43RSQ9/6Th1Ze9ODHMH
1Ow/gANoSEBLB/SLSjfLMlWxzSx5vhnlOeJXy+vVwPXDGE6XY4+UvOSXGqCwkS2iusUpDmfbHfis
612yVrFmwDiyPEIDFhvGxzxfjhnkvpECGQvz7IstRp94e9GGE6nWReS4wNrpaFXeO55PjK3VzQp3
SKApzJFTsU7Ik7Ds1uWIVAqr2Sr147pmbZkCGKWM5qM02jnpZ7JXNcL+YzMqB2MAyMFnOKddiSHU
WD6x/M74XmAvMPz/FdSaQUprlZTIvUlm3t8sEe3LiPjjM68pz0hiuW4Oq/d8dTYbyEJDWbnyfLE/
FCAXBpB7Qcb+Zufh33IIPV5/uKxDWmOzlzYxkcGvFJsALPyz42fWEdgKs0EaXQ3Lt64QdgveAFWw
+Q/ulUDQGLBGNRzgkfIQY095JcMiXSFzNbAJRJcQra9kjBlAvEp//XjIoB7OIKdRAI9XjBKd2cOd
5EuO5+Fgy/4VoceplKffKowXSqT1p0gaOO9Xvr/sUw8IuCsfDNFTtKL9dpytl1C05/if+It70+Oq
lFdkgFwTjUwYgyHRuV9zAHP0+23drZdu59Lak79j1wjQjWBXHrZRZEXKHyAZKAq5SqTb6mxeU/eF
tCDm5V5GLDCqMPh4mrQsTgtcF+CB5rXfPgnXIr0FBDOupKj0VDtUxBWdHa9PvnpIPcjBTbcvSVYR
rORcyZx29Tzrn/2bk1DasBOtD90yRRmObW4/gfAd0oifSIpEd84uRoGrbEYCWgLcGAyAkJ3oc/NU
dVbOVUlicDFhWdpgHXIWgdxDvncG2HsBWQLYpAilKBKsZNGLF0HPcw5qup8b4jTj9+3ieU5EvcfU
t1WNNWE54FSqn4MpWR3thftZBm7t7Jk/fWJSLMMyJ8Nc7hIQsI3XjTsnONLPGJWejyR2p2sp68or
gI2XJ/9gwdJcm6TrM5KU45zSIEw2eXphyapI10z/5wd8cF9yVuhFWS2zynDAivSajSOz0EsXb/hB
Ru7jYw117HCFww/noKP/v9naEpYpguGakaLttjsuoj1og1JHj4IzXpVNwSozrcLZfkZ/A7o31ezu
oqK4B2r3OV+Wyx7TtLT0PVZz1IBExq0qhJjEu/LD6neLVSR1H1UeDMI3DtePUkO5QjDAJnB3z5Qb
OzL9OTxYWU8QzC/kKdUnZ/DZSVP08Ljf6qm35pTXSB2ubfrVb8kOfzhOf7lQc7PJnn+H2qlrFfTB
0DTkNuGmSO1CJpat9hf6hk4VuuHvAhxc9W7IW6n5dSt3juJJst/03t7OAB0te6cw9cimtru0GqC5
YSLYnWjGbRIECDSb0jEC9e33PUKmrx+CYmFN3iaaK77Dtof664SAWh3kJGwt1qm5mZX8mYq7T+Ft
BEPSTqGzHY5Pc5NOT9U/jl/0jj93nWme5flLJHhHdN5y83M8gIDmv6ZZH3pdzu29wxFr3a5UYJhN
rRUytS8nRMuLlAIbPfG+038wp8lOl2J5BiF1DQflFGWPdSEcXrj0ITdIoQb9JuEEcl64Kiy6n4lt
Ug5KtfA50VhbkwAFBJ86EKRXIJ11OKbX9G9JEcr1L2a6FhviLqXnn/K8ZYqT3RGj84LKuTpTlNLy
9DopCEhuLwdl8z9HBUZ0J9NRLES4CoumcJA4FRbCN5HxKCOkcqjiwn4iz6/dxXIHL6HvQ62CN/Gf
tL6+WIs/HY46CYeqftiu1NQEhMLlTLKBXqyvZZlFl/jdLbiv9CbUvIk36U1yRB+QbQIV2J9ngiiN
sctq1ZSyeALio+0povy8zPD08MEE8vAje59rU5CE0jI3kk50RoIutf1pK1RhTAefxBlwVnC6pM9d
as/7/OKrloyKl+nTtaunKXBLpUxdvIKAlgt/ZH6Z6LbFCvDz/YM5tx9DKovn6wezG4Bp78A0l07V
CJPvbTdm13kZtgG24cKnyjO6SGvbFw0nB/ltUXKTY8JiTIsgTDOC4DRqCAwwdISuHQkMS7AYgHea
MdGaGisGXgyrSZbnR6caCunTa5GeJwui9CjD3b6EKMKVS+yWuZzjAyoMCy3dtOM3PH8UoXLnJChM
nESVJpNlzdWRCdEdxXLLAlkSFWIQJAFHeAwBARl6kjj1h5Sa/QSFnpxFkhDiFEzHknWzYJsmPeZ8
4qN33R2q6yEsa8x6rrwxO/rm3rCztxz2+4dFATmytbDmctDUgQpCDoP5fpnGCDEXDXNRfNj+4v+Z
lOpinS948Vq7G7dcr82stLTAeTyeh7FjFwrWxXQ+OjC+oXCRUSYykmTX0knYiLD6ZziBDzApS1MO
9ASag/mkFfrT/gcXB417bXIHkNFkO1Ptcc8/Jsrql81K2E3g/DToHXXboFwP0acXIYapGwggDzD7
XqWooZWfWnmp2KRmSp6l0Wl5Sxqe+GQquoTWBQhDAWNQ3vKHBj0tjkVJ48DMzbOyRRGSuralCIdc
Havx1GctZsRZXInn1zGmuIQ4t4HjpKjWfwTPRhkC3ys3COnXiy0ccescS0HMidb65YATetT5Fa5G
rzlyUZivo6DhZyHOtswOw7jbPxEIWzlPY9iSQRQXPgvDSVHO+3Gov7Bwe9rQBDdQ17CwUj7L2w5a
tkRhVtmcvEbVR4v53C5iBfkPg3K2LSz7oF42fmPQPTKA+moNE0ufOb2fNykIL+53emWXGK/qkOKk
XQegSBdI4aKbwSwswIdCHR0toLorNRjNtN7bxwbYiEkSpvzWqQ/lmtawrqirIObUqzrHnOc0eE+D
rf/nVBQlEb4IvVzhZR0Mbz/lqy9saz8yXpENdSqrop9wEAV0KuHs0ahInJ49iCBPt51PaGM+yMLG
cK/lcmLiFCCJLBX7E0Rb0TSOAvLtf+MuyyjpEPpmjg9bCtz+mSMtwHOt418fYOj5/m/0ae9ptNcZ
KmG7AqUB25ttGFODwGLcKB65dYLm9x0lBc+zJkbpnLCVAVpuI/zqC9fWF8ltVHh7EMVau5CTaVLN
Vmz9Ll7e4Bg4VvLNg8Zt45T8YlrC14lvSNLzZxG1yxRx9OJy+FaZIDVxESAc3GCDeJF5vwNgnZ93
z+chnM/fd/6TLpE16+mIYPOGtg6pZlR1zPWp3xcdTStcdVXZGZ/9754AAxCQDzjpyvEsQRM611pR
6qp9zfYIExZIw2VuPdgHI5M6UXhg8ULyeYZVQ/Ct0yudHQvZqsea3UohgFHbPGb+oEECnddHOB5j
eul70a4syx8uFNEDWKzyPvZi2XPcZKiGw/+l4jJaXhnnPbTVIWt4rh5uKc3zMK0Wl2WhwhxvXcix
ycLsWHRyYp4hg1iCuQbnz5cOGnb0RD1GxccX7t6TCG5cHr7voE2UeznAPTs2oLNHnAekE2fFy31t
A/LuXxuf0rnMDJIdsS4Q30PGo39b+ad/MdOLpQTfgI/5EHt1wVAQf3ipAyLQaQadkfNFgBP+56rs
DAsLEcnr++myrMipqs5a0GB11BdIiQltEpi18Bv9gSY0bZEHIYwOTUD1VKgmPdyYF9o5V/9DdHLm
XK65vr7RtqTxOijnMcOC9Z182o7E+e1AISo7U/0yShhk7qjS5OpBxwwxxq8qlBLQa4HSFbb47edr
B90xXS86PGPvQfWf2FxAJW+CK1jhu8a5JPDM2S9c4RoaKO256FoeRtSq/l1lC3HcdYo5w28ZwQHH
EsYq21XXD/gDdMLGq/rNmnYZL97Nn1fy9Z3Or7v9IBOnUTkP+E88nN4kFTdeJHH3mXug5+46ivqC
58vMl/8bGto49cfwrZNxYdFbSfe13+jNpuS8b9hhglMk0A11GmTI797K06h8dkxr5gxCWb6m2piU
dB++PcHdQaJ9Wz4dicj8vWz5kYNRBl9834abiP1+z8v1YWPt2p6Q89D0zYx4CMT/ihfcWUZwhg5a
FvaRJY0Mr9sm6yOwTATk+UFek/+x5z7Lvry2F3bcxBq7p6qgbrt0zwzyevs/NWYmJa8cFROpX8Ae
k0JlzJoMlWXWPADTXP6ZeCn/FoTeXzlChxtocbszj9aB0tvmLCvhwmd3I1jelmoQwwee/CtiG5WS
B2ndkwqS1x5uE7HRjH5e4XX76czfjTDlbSCVDcJwh74lk5NCdadX8DXEundznkPxgpP0LM22b20u
YUTuXKaAPPpGGYrXaaYWwwO9gjmzWx9/hG8Ms/tTUofZUDE5J2G79VJYIEC6G1uvWraBVnx5kumI
kXzTP3ZEQyPWSXu2hobxeaKqTRfbJq6Njxie2Hhgfy9T3TnlBbcz4GLree/yXdbZ94KFjJkhuh0g
Yx7FHNitWWRFCKGKao0kfdLPnZLkz1WOfkl07ZPCHkZFBO6lWYjPXTD4XDEjVpA3thcW50ZVEVdr
tatCkCP1blKAl6B3Gws+6NJt5PoFzTJwWJdaRcJNdsmK9+TQZtMvB4BcVL1xpln66hPKKAYmz2Mi
yt7DHX74IOxtVa57Gy7o5aNrcPp9GSkSjUlHM1iPmFx69dTXFoDB1IEhsp3Y2+2WQLdCO1EhiUEh
Osix4FhoHPiLmMW0SEXxR7ibqGUSe/JB5UYpIZwsFRfpFgmhWc3DX5znXG7yTVj4ynljjBlUIuWs
K3rDWq1Pa4DbnGISSyznolXAKTdoy+CPZ5OI6559ywiFN623oMNk7Km5p8XMmK5zZ4Srk8Fmi378
3v24K8kC3Ky21LB4hUkIif0t/6TQhj92S1tlv+woMybbCi+TrzXkA/DRiSAiYM3IWXh91cHUW9k8
wscqixcobDENoBcoZeVPdj2AFYw9hubDJ0yGAWROjatsB4rPvmoVPpxVBe1S4ARKu0JAfSjHoUlX
BhNPF3ihvRIp+qYZtvfqeszD2x/9UG1n+aCFR1iWoNhWeXSB48+zPpF/9XMPUt2/JwC2ToBnLGPY
LjJmF42ofmsZ0wg/uuyLjQshLjIEtUnd8V2t1PuYgTzUJYAK3mCqArB1g3aTN6YGMC4CNtFG5c1z
ANGAeeDziGgjpAa4/pJT30VADHZnR5DWjL+G/e4iIKJFLtw1BW1ZnitxDIt04P+xZgIX97ddb2Fo
cY42lHz7wy20KqgAn/NFvvA1VL3KLaFSypwJ//vncMLHNnyyzkokCq5YAAn+/VdnXQcMJajwvTUf
QXuyltiVqm0Gu6s5TIEW6Jy4LpZ7+2SzX/Bg4nx25qZ21kqu5+V05ui/sm/1ec2lOSPEmA5d/Ds9
pMuL/QxWkgagl1rim8A+8W2WhGpp0GfP7cUaqW+UP1duS96yBUlmhOIXfgslZqv/9G1klq8qWCwz
3xp8iMkAPtJe6/5KhAPY1AMorDPyAw1kO12a5mlb0Feg/ugP+fseD+UBLaGP9AVnmmxdbNW8uCGl
VRUK9U7oSpEhk4fmBZmmtun6+PXJavAoinlhMyEo/vt6JD+oHG76sBlGdnG2MJ/CkxMc9UN6xDlP
5y/kh6sg2gfXRQfGrrBx7bdYl+M8TdHK4sciyicO/xuR8zWS+Iewxwd1N3haj8q9MJBX0fuACC8H
i0y+5YI5e0JWdjR/dg7l3OCX0psystkbXYjkahy1fNPLUYgBJ6G3NLwYI/X1gpLEM1f+0ejNCCjv
KR/+L/e4Z2igFkF3YOKw9+uCA7lYCDQEjHAhXSPczgRMVjZNFovYobZESp7eHpGiErCM0R0f0YCJ
1iKUTA4NjE+zp8AmN3eNTy9p2S6AuAo7+XV2dEhVe/Ovdu3KjqDGS3iFzYP/aBsl/93yY/CD7SY0
9psIWzd6fWgJclHin5lphOvxEqP5uIf6Lwp5PkwYsrsyky34VHl0pvEN6oRHfMmH8K1UL46TkT/e
Ksj78u55J71jtd9P4H9ECial+2nxTXFeF30AXOt9qSDLfNElrHtvL22fUWN4xYunszw952E5VS8b
y2qia1jAoSx6jIC3qivtVWVTYECWBTJHe4Hbc9XCpLeYsR+XGvydDqeKVEVXLHOfaWQ8ATv4lQCL
IzL4LXFdRjzvNASfO4JvHbssXce0ufmx8KBwMYPEFYHo7iSIMEXPL1Cj2GVtfS/O6gS3DJfdXeLw
KpfSmxEUvO1HA+gg4D316IonMWrc4NYSi0WB2LSezXkQZau8mtl9OvSo5pGoS6e5Tp34H4WJ5Jg4
QT7l6OEtp3oIeScXKfQK8jjL3Bh2bHidrbz+0d7uhAoO5w54LSNzSqTSZdxdy7nthI/oFDiVYpQ2
mXjMrPxiuV7f4AFg+wMumLussuiYcfu62dWiuvbmqOZO65xgyeLiQN7WvwoIvy5D4kLkN9SWg9JD
sXBIbt7LG6PFDZR0kKDQyka1uu2rQZ6tR5fxiurdoc6oO+cE9Fsk5ULIVSXqzl93CPb3CPVR4+rK
Xlj0hvSOLTOlOROcgpxr9Np8kfqfsgn5Kss4BlbIPx8XXNjv005/aCjVCd0iFSZLt0pYj5KcHbAQ
S9C2j7PDcPFY4NVh6T2g1w0gzhLB7k2zgsLRIzVdR3iS45IScVSV4wD6Hz0/jNbZHm9qyMTNzgI5
cNnloitZJD0G+RKnI9kDZH39lx6/nSZh+Va+ZQ1Plnfk2RVgUgJ/1OXGen5Qbptj8i3rEIh2VIsx
46tMfGDRR9zlz81SB5vufaJpHplqGzIuFJE3t6KVa6kD6+dn8lwatnvIWHK5pHWlW0/tmboIhBrc
/Ue6nMKH0cOZlZcoGEo0ouRYU+zOclc/lBWcCGD9wYO9dklubW19S+0KStAH8wJwbbireA0AG0tx
PlSEoKbe5dDSJgm09gRAxf08pZHQV2UaTCItH1BLpLTp7VC/p/VRMec1Kma+iy0iObEQ9v0sczWh
yMrV9qVwjzlMjjktOLZ9xFmJbeIXrq8fNMstbTnwrmwKVFM3Y4gMuQQoRkAKMzMdj583x94raSjH
o7dDPzc4y6Ba4X7mVHOu7hvb5jMChM9a0+Mq57TH9S6mOq1J4OzuKphWBd0ARFbf/cerh0aK9rrl
mCU0epR7UlV1OTK4q7oWTUtR1pkNxI05kn6iPXcH/mZ3yO8QBktP7reBKAvzzkzPTeyQ105cSsMO
wOlsMgOX7/ZN+Z11Ctumjo2N4r6NMncL+fqPVL9vqIy7AJfGkVg456G08dd27GrX80jepB2mN+Be
SyKpry9pGWI1NcOejSHjma1/xH659YPnyoKlUBTDQalhH5DxCfcagYw/sWB9+0V6WFQ/3xmE+LNX
/Qe2jf8vJyqPj04FZXoQCbMtH4WDDPJWcCnpcUrT18MPtCnLLecajO0LcimozbOuiCJRLdspDY2y
lXnVVznUxEN1aKpbCl+pRLMpA0hw8TbBUWt2OWlu9fxr139CgC33Oob1rC6bzkhfsdT3wWVMGist
4yZNTsgZrbiiYbJ8godeI7d0FlHA6igrymjb1dnlOysfKrb/KjKPu85mpl/ijonmL54BTszhfZIo
A5o/XfHk1mDSSg4TNPl5aURA/ArAiR7QVf3jVrIwO8iPpd9F79h4y0OKVDhjGvQWwUOjNC4FTMFr
7dRrmSPzaZ8x9l+W2Ro51hKG7jBtRBRexYImqnh59uR+z7CPseQgMnVF0Qc7OuM/xi1lhOFXuCmc
isNvuPJa0mXFOKgBrCgunA9Z8MU5azfGNmqUhT6DiRY73pzCRb5y0EiJz80UkI+HUgW1fpt5LWau
xGpyhP/3FVjzn63SXiFZ+EsvWuC6mLn1rjvdKSieDmdXTTMK09551q2eQGcY8RR4XqZ8lTVfkmjQ
5LQe+4SxLYyjAgwdO9NJWN//Htg6yk4PV1WH9zjaMKHbtZE9E2h2FEg7F0a/oKd1guKxgacC3cIy
boI7rrU1R0+z6YMP2nGQCZjJjeRnBmhN6kaFHUNBt7YabexaLDkzHgtoYr85r8+FJO19rzA5E0ix
3RZxc87V7waN/7Uwhb66Dl5qJqUmlJ1bpo75CXsf7+Om3f+XcZ32C57T7KyZzFISfbwvNLg2PL8g
/4NGi8y9nBZb/z3XLDdoFB7DexVxc+mBEdo2DiHtrPXpZBhnDovvIuX0g5Lj1sIPBk482soiA+I2
GE+b86A67nfEyA30XuMXSQaGhm82eLFTZXJ6/F2wA2UnfWLcLHzORlKVj5kTuz4T4InCcnONQD65
OGFOrRrRripum0ivDpxOCJKZQp0wvLSi4WSpCaHREpr2NXTzRxvh9f/eAxjrNmKHavaxDRrqn04D
PKc9DcmA0XltEcSk66OGMakAcuucbAB6Vrc56tbN1j0+aOHClBZf9vHq7Vu0ZVOIt0mhOH2QXzg9
hv9yjC9bFMJbRrV6Oxr3rutFkmWyw+rL+FWpzGTsM9MyAIfMaQUeA7WPHCy73kTxs2ARZPAVkSg5
YCeJSKUWI1qVTl3wFTO4pZt48HZ0bazPwfXnXYb9aeqmGmAxOShPbbmXcHTzRt6pbuG1Y5EWzXHX
KCfT4/sPH2eJ4j9L8pud4rJoXrpAwJou+V7TIEyBxCTNAEaZ9QIVW5O8Se91VxpLa197UqEYIW2t
0ioCbMnibAVlM/oTOc3UnGyTJb/OXFrxDwbXXdL48X0wzr+C9JFtcbOsjPpAv9otIJV+r0qxpQsA
H8iVCxGy1FYpBPtBuTfBRH+k2WX4iPnrLj/v4fQ8UzqazSye4XrTu0+bE4wIfaZgoZD0Noit7nOQ
64W/uhg7SF+lxgrWi4TKBEt7cCal+lpqsgm5LPOewO7pc6SSHOns0RyEIUzM2C2lacbplXdZdLux
G0H3w4TWBqMC6DQNOmyL9nv3iQKubEzvea/wpZLRA3UFrLPHg6RcJxc1oyyYpUXoqOlQa0QThmKo
y3iFYvebp75FYkC9lFpJEvABJOD42ZcwAGfsN+qa7wQ8IDaRkV1/5kgsYVqmJTAZ4mB0ZmtspPRI
0zp4I5Xe83zxdddLv4hMQCPzkTSlGHvKzeYlpWGUPZsiXAJ0l6ScTIUsqn/d7YL9P7aOHSe+HCXu
Fl61QduBfcuPDKGv3qZSvrpDSgrYNaMdYlC20g3ghNuF21Gpu2yQVX+Hs0TGE8PLU4q4awVj7wW2
dBSwmS2FlfFGgMvUOSIKfq4nNZr/TplVls51BQcXGzkayMnbAIkHu83olujQf9PQ/S/F6vy1RJUC
x1XvMn1RcSPp+nENIjdJHPFOYpNTg462MEAnqEdc8KsXrGOpAXYQ97bR3e0quJL7s4aPo6hHIYo2
NmPW8V68Xmxqhd4C8ModIo94VGQv9HXS8P2p7JaEzrYh2dBBK/PzV2hjbOoVLMu8s6+TxSBjGwRL
UHHRBRGjvdWMB+8r0jmqXKk3x1C5suBmul6iGl95SaaC4XvOZKDR7LL0HbsWXkAnb1A95kjW1npS
acB3Gg/F77ju65PrcdP/BP6K56jTp5E9UjMnEy11J0htq+/uW/b0HhWnPDp1W27NCiznq4LaZ6rv
KKKx2eYy9jNqOaR6mi2tyM4T9P2+qg2CAeX6r8mQRX3pyMfs4WtTDM7i0CoN1OVvXCEPYt4zc8tU
4QVf8H/PIsIt8pd/4lxd/5YZ6RkOknNxgaNddguNDtD1ZUQ4hnK/bZIRdvtvUcrU7h1l2mOOX77N
A8sFn5eegbdoqQ121YKWLxuUj0IPMX9y4JuZBzWI/P35thxhHm+b+L9gZPpHSjQsxaqIpH6hIzCR
GAE8V4jvA1Gtmfthp+63UN4+7F5B441g2NIElbAsajtxbOXaZotmsQo225p7H2HJTm3nuhv25odR
ArLx7NWOYUm6msYJTcTR/EHY9MOly/8+2Fjns813Wdx+kQdIdcAmVnuqT46SvxLKD+fKvoeQFzTv
0Fd0PV7IVm9fI3LKag6DEy3/i0/k/Z+9wGouggKejxEXbYJikTUi6wDsszj8dzfZ7m31fGrKYBjm
tShdcQRUJDdHYXQM4LfHOjTWShIJb9zI8TtEWFncb/tV8XLmPTkVxnXHZsfB7bgZ0EHb7HZghWlT
NfwPQLPSR50vVntmjsYuTpISb/qX3a2/mm6NR4JUehtYJhpqxxa61bvkbPB+mbSe4YEa2I9IlhBn
+9opPDi4l/RAx0cAGtYZlKLflzP/l3ZFGUm0owdEHYfcArVmQiLx/F2USGpAxGgPAU8xXAAIh4v2
M/izP1wGFJRF4jCOQ4r4g0VgieZDY7pbpZ5qw8KGo86mPG4kDtBtNGqeR14WCIXukwdEhyGAwp1F
6nAV8WF3q34c653bT4TlcmHZGSqL+Fl/yo/799bARH0qjXQhzZaOxxMdZkjridVrC3vhnUbgmw8u
Yb/zGv6bmMQ+TEatH0bGynO6PKYRj6KiPQ0t5oeBEDTaCAXxbjSZZddSl3qS9nJCIwa7B9QIGAIh
XtixWx6H0LvR4kVvAmtez2HRD0Jvm39aENatemKkPHuWeWUtG1nJ1qjH25MCxscrAfRpWLV3WDKD
7mIhLNOJ1yVrgU/ByGJSetXkE1OHizDZIgti2zIUXGv1oI3WE4DVii2UM9LUwBS3nkLsC1cXq2K3
dVNLmZV9PeCxLgRgjXFEpsZlZk2chm0AsWJm4496oNVGy7+mINBxDp270ttk35hKKZileWadjUxR
54gLcS+Z9wXxBGkPuzXjeZLtJ0De/QT46ZhDCRe25otWbLUMzS8qZgpeCjyUf4lzMokWn8cB0ccc
PD7zSR0dcC3lwIZ0EKhvfZGnO94iaMPruVrFdA7mUx5oLz9e6yNf70hp87fq4jZCwHW758x2Ddho
Qn7pu5+QXxXmJZdjBauvZQtIu967NJSP7aBq0crGaihnxB9k2Fx08r3TgyiJk0wPKEtBqEpCMj2S
9fmXAK73fveJU+P/wGCqBl/TONdHsk3lg8kgaon7GXn1aDRw3+A9V732XQ5c5Z1QR2hXLMOAmbjC
AuAKzhCeKzW3lb8+CIbHdUzCcR4UUWjxyq0ajvrbnHDzEKnl59Il4erAufMnYCUTb9h6dUSvyKo7
tBZkU0s1EQEwDRj1SFQlGo0F+AdsRlLgJOGcYQ82ODceBHhl/6VCwTSG6TLrddR/8b45xjfu+2Zm
Q0wsXkYjKqja15wW0O9Sx/1XltCFP0UitqHJO5ioGa2HFxTn4cQGnwzI3Hpagb7O0xyvMR+jzre6
4On0HLBwBugrJIaLUF7OnUxQQavr8RfwCgpRuy0cUDBMo+oQEXIr7B0XSj/eLm0GVLGZQqh1i67J
Lu9gsdnuY0XjR/fbvt0eZRBssOY2BGyNCe89joOS9D2X8Ei1DuHm0Ku8Ymsq4DuP6TX6jcpVc4nS
Qkj0/KGqFEaeEJOE92kP3SPx1hYCJQB5D497IoWfVbknrTzz5qhSP3Tk+RuqVwEStQMbDkxPT9IZ
fopSwf3tU1QAJtdmn84ahKG4X/vk4iDALdj3pU/O1IIl51F5OpGQC1X60RFGa+I8z3qBZKMThD6Y
wpC6WZAFhP5GAQK6S3kSS556wyAhsazrHpy6+/AtbkbkoXFm7L8JaFvgyGwiyYTNuqkLjhjosuYh
A4+bSNJh4bEKrPeb4hdILY5Rl1cLGSBGftTJWnKzq6YaPwBXOTThVY4ZrK2X10wZh1YRUxubL2oI
XTnssD8uk4jae156sZxR1PCUHV+WmZVaoruvQ8UQJDtGUCHOLCRMM8zQ5ZY1CVgpOBKnm8JowIyF
wGBKGxS9vNumBgE9ohLZ4Qs7ENXV7pD8tdvspYq47JVQhCCnJ9gEWRYNAGxcShMkAnlG/EFMSMzZ
StfzmMbKo9QBMY/Kf5VV4xl39in/1hwgtIZFbQ0DRkZHWSxyDcEuygj41uIzgb0Zs243aCtMthRh
h7AWLupI4xW3oLcqbj+RCLOS7okuyy4TWJxd3DjFsuu1uIv/j6QF9IBaJfO7cjuDMbepcWieKvdz
n0fI22CTBtUKGHtGjwP5MeUYbz/UJw51EGMDBICJudtgPornniRxd1m+ZD5gjr/O/bzj7T8eUqMW
NmIEZIZx6xkZwRQjVMeFNCMIcv1pvfs8Bi9F9SKUy+T9x/6CAQgn4Aenk++YtPV0cQPh2ljuq7E4
JVovWSzYP/L4MgHq2PW3kaoBhnzummIseyotSM1r6BRE2BLJaGnDg4cmc7dhlaWJGP5u4ZScuOwn
VsPeRnCNIHKm1GdfUXACUOeRWBeBt+mxKnFRgWMkwP4rFtG+/qqVfL+n11dzToKIqHbo967BY2/3
unWFQKhHqm5mBQYpqwlYuEOoT0idLIlsoItYIM566tmNTsJYj+GEeSDoMjgFCsY8RbLqbS5G6K63
fvsOqjwx0cWi8b0Hqtud8OfOdjuq4RAZz2f8z49yy2R2DXH1bwuY3SsqAnZcXEVKKXrD/62if8Ak
rAiCQ8DXOZGaI5pzwoxlQwbEfK9V/z8xoG1PpDZrAQiiwwf2wriauvxLztlgHZqHTpL0ymej69GG
iGPa0wkmGW0QWA1puAQIRYhQGl1WTiueZ4sENi74eM7gI3O0us9xVmxG/sXWBp1sJx6cWlNzFNZe
H9I+7X6kFueaRrM9T/RkOqLMZWxMlGiXQL8VSe4/fbwE1EJmWD1fwHwnWtaK98/YKbT9DH8L/JP1
kV5MnbxSeTegJh18D+RNjBTA17DP+++HRyuzbiXhGTDkJeU0gS2u9pStMU/sLsEoIH+dPnJiOI+P
hRBG8PAWkCtpa8KErrXXJOeZ+CPQ0hGPEMYHJ2km6O+uyYKiFEKccpa70Ib1JBNadqcZUoiipWQP
DnLgYJw/Idlx2fyC8yz+FuvoKewaEoSFV5S4kkae1GZpSm10vVITOyqxQqNdxHwyNZtIyzEGSFD7
blPKEDRMJxoBlOKeD+iYjBkR+tJomvGOgYNjgfm13Pw3pLcvhAcgmA0TmiyH+l1Neua0q9eGnTLp
pCoxguuwulzkwBWG8JhT8shDjPt5EbP0FfjMrdnhfA+DMk9zz4z69duV3z6354dRm5hCVcpt1il/
v0/KYYPPJ1VOwwaJyaNfUv5svSbHNfMIeVcU7InQsL2YFfp2FolG/AkZnLsUWeMye8gp4+fj8hut
BxYwSIadl8Q/b7ccASwfnjXKDSA1sj2xOl0010xdl44bIoaN7pgIUH4wpg31/ye/FQQkGAfPtseK
+RvruPDPagW6zrWwwqfsst0wlH6C/mzrydp7tzzvz+50D/p0rcfFOgjnKpcDTwBAbHljj9Cf6fLl
VH8um6Mve2RsiV4/o8lbZaQTzsN5eK7EU4GPWZSbuwIe3T4UnHiJ3kcQoAq+nRSIy6I7Ae5YdbtN
ZztgfeN/HIiiy2YkGGlGXp2hSF6OiPBOUNtA4W2i2eiz7H2H9zgYk40MmwRIyJzmDexpbozXdilD
kDIJQq05jbiWuqbd2/50h7DzjQm3G79ICf19M6qEgC/Wx1NfysJOOuXE9CWWuGjZ9/KEbsuuC3Dy
oPlkRVWIRSSCnYpIdtgxUXqg4X7l90293uxbeqStFd/uEL6VttUemfmbs+sP+iWPPfgDbmo9LBoD
5kebqnJTpqsMIUbTHn/vN36HQ4VEpQrXJMeNmxpMWfMvesveaN1dCPd8PmXNUCuUu5qEXOa40wqu
4RmrHcwbidbxpC9zyk97CoDs/+ofyW7ER0We8qFLlVeI1Zmf8z1VL1isKbMrV+DUQNSkt5DuAlTD
i2fpvpqSequgkqPNKM03cBp1AW6wp1jYFgnWhNGqx2aSVTenIQtNHsQzb8K6mmoUHEX1I7NY48Vf
/ze1h3KGrPJCCGFPpMxn+TQ/p0TZmfl400Bvp5H2XoRr+1eT0c1AJt+q3hBUmJhu0k7eI/Z+e0Rg
LEB2IUDFqceraOA03KVoxiR8mRcRhLk5r0HUlKTjHEsHrcIrXX9Fq24qRbEP5Uxnetb+4/U0BJP1
p2Q3/I506lrc65hCuOYG+OngVVQHXLBhKJD6rfTIeg8gx5mvAdex3Gy4EhWUO3ggqmF8gwWAJM2V
xJLzUW+rOWba2fWeNOaErnpyLQO34zEtE002PT+w2vstmc5BdKqmbc83T0KCJfcldUkPEj8ierxt
Ekw8yfE8nAooPcYWnystPX3ez247gdaPz+FeGVth8eM1LvfpWOCaXMD0BzeuyNU7tLJQbe8ABaaP
11PJb0wYEwFEjJQuuPfuU2SbBP/xbWcDYyYRMakWoaCOtH2OWZGIV0Oa6otAj041Ykf7eJmjbOg+
eQ82fCslPiWinuuycdWm8AE6MloRUkyY3r+9uSmv3qRV40rTiLPAc/pMcTtKCo+fSbkHJGhgHcMt
ocnVUcg0VKnx4/4cJghElUYiyR6UWLdZ8iIAyB8KkQ9QcweJqDr99EenpyPtwSrMQhPCVHf7HnZy
fryXCkhARAD/5rNYjxU1E0LxBwOjdG42I/IX2GQvBx/19yry7lWtOW5fSJwAEOuO4UaMNvAEmzYe
rWmWJV0EwMuWkqkDQbg7c/7jAWMcTs/2Dy9DcyCx8VZgmfYoHqHTjkAxNQO5zLgb+STqUdygwyBR
hFM61D+UM1Lq8tR29a0n5g1VIoaJjcvm+u781szBMZrhV+0UltikY8eiG+OYi5cngQUDdRpV/ieb
fTPCah9UhA3HCslvYJfn6HEF4LFb2Cv4lUfE9LtHLgssrD31KpPQzTSov/jSly3xde540lmW2kZq
BRX/GZJ/MT2uHwM7DFus8jbZEdsgIkZozwpsZfMPITEvcHSkXUEQO9aO6Y7vmvRIplss5FYWeNcv
gU/fTkYoLEiA6mGFhxktOUuJf5K6wJscy+Y1i484ve3v5kJ3FvYoWO9Hv7A9pr6q+27FUUNMOhCG
QDPtauUcR3ELVRpgcjeYNVxZs3osqwt7z2izcozwqGzs5Ezac0blWpRUIxHILyXLRlss6EK7Pe20
SMGCseT8bFIDVLFNwFLzKsGF3Vg+L1PKLLDXEuW+Xf0fFcWTgPhUKzVLfb2axavLLsJwsJyUwma4
m4DLg5IxWTIlNYEuo9QB6hnSzFyUetMHvUBnsImry6+5ZTJT3OY5GFliaYEIm62q+m5I/4LRhZ60
zNz5g01ORnqbzAWHCBoHmdG7JpCLtEwKiM8PM8LrJAkTy3N4w2kMP7TXnvvjyXzQeRzmCMo9j3aN
O/H9eL6XzYkCpbyndLRu2YuoEFwhN2rPyq12FXKTobCH1ATkIphlKhLt3FvDN0KNLMYiFMVcfKyT
1z3O+5SlTSoD5wy0PZdc5+pkVqhr3xbmTCZ5Pn4lKESLIsZVd62NdsXf+npy5VfWHq3cxcQCDeAC
pyEMtzTEe7iFU1rK8MXWuNdD0Toxn2qHUiCdP1ex5xg1bERorkieVOFPw+KWaRyRjD/1+MccuB5o
UAHZwfyz2nhysHYrKok8ayCwxVdFa0k9i00N6SMvE/jOtz6Gim1bDHBycrh9pmqjEMGdhunQ/rVw
s7C26//guaCKCjROXTQH/8HDPTsEYbJ3f1BRlSmDtjyiJbvFIElss0Htilre52EoFoNRCe/kST0k
mYVLQ9izstBOnMPwxoZs1VmOZ/XQ5+eEBiaYDziJWe+FeWRgHpC6gV6or7hJdnmkhTd5hq1wgKAs
HZjbStL+3hGw0fkbW+ipzFpBAFZ5NO/9NAVEWxPZLCfWJsug6ux4KjlJGQsTbcH4kAY4Ny7QgaAi
6G0iaBerN4fmAUHNcc6n0IzZg1uteYHooqMSyayNol33/n1B2HYugj8AHcPk8mKBtOAmrjaY/eaz
3yAad1KLh+16Vf5qeRbftHcDK9uOD47+9x1vlGZYmfWlbt30Zmf3boHdqYzyBGZZJJUBSHHu/w4z
R14XWn3MUBgGiOaI4INqoGYQxxLUgLQULG3in/wckSO/K+o5I6BXQonXIwme0LVebcVdriRntEma
Oufx84N6T86ZyREDFv5N62+NftSrteQm6fdkWrFkOKx/ChGZCieIhpGW/62rGONOE7ZvtqZPgHPm
KVpna71dHtgC/3YsNvEH5LrA6+HLk0YAij3zoEe7BpMKNdrhq0ylCU3Pd1GXN64ve0y8pAAFehc2
3tTh9s9m88bF7X/hkklBWkfnbwMJqF5u6f8554GAs51QhRTYiOmooFxX4E4BHSwZTHbA5faRDs+j
O4LSMJ7AmlSsS/7eMc1atJqL7pbWwxoSnJbT9xPBUXjTbXU4Ymh+QTQ0Jv/MNL3iy6krXZIAbRT6
Wtq9P2HV1ms7/4oeTZZz8k8GDviRcX5UMh/jYrNxIkB5lBnw5A9Ao+Gu3nVflFMNf07Y0zUvHDAP
9DXAKlJQ5yWdZZbbiU0WluFaHKnzACb3G5EOKTRxWwDW6jleGrkUtUjOhfUdyIelYLy1XBpbCrQi
O+RyXOeInT+FVylRXcuC9MOK9CK8lX9lcfZuq3b8ZkBx5w39NCbhcjL0827gUqQwJqXXR7XFU7fT
7/NBasPKgPdxjAt5GA5bC/Su+eCIMKe+ozMaGL4Dd9gQqFeckFfnuQEO2Ko3jSos9RptYf03MXiu
EEBCLdJRQGc9iW2HyFi4+tN8NvUi5UdXgoQLHCAWkT2hQDnicznd49xcyO/TBkes6jsox3Vxv+Pg
xcMQ+aY40VTTwF+r/J1DLqTIJJL9leCzsWD+reQ7J2BFR+H4zYEjchhnWvJFi7J5/hQxvdezWQzk
gl4qKT4dq27+EPVIOBxuB/x5PjzD40T6BipQQ3PMdyZ3mtpeXMO9M2KMmpROYh7Hi9xUZ/Pdp82A
wysxt4GIw9D1QYAm9HO0MCZVOJWapl7q7bFU3PFRLatKaP+79hrTIfoxrK2wlzeDiNwwdAAzMfEO
U0FdLNuT/Fo/jnLQ1xCKcsAqnjAOhmwhYqGfpatlCDRvuJxPxLvDNUt01lORk5VvskhR6G6nITmE
StS8IqLHRsUj+8n6ZZSmJb4LPPWxg2lk1CDHgBRkwbQyrZhHo7JBtNT8O1roXLVq4lkg3lnz+hni
9CC7LfWdNo8rEGY6hT+kEME6AXy+5JKsi5uNfe++/g82kCWE5S36qRPiAlkXww0veD27W7gHp1zj
wnu5Mh5Y7ysEHHANPZVsbXwqKeeKWODuB+3TUlRVRQHLN5n9KSR01Rqpu94f8wXB7n/UEgDEKVpl
oiH3d+YD+rDOcuGf4hUumQ9RGOUrWzKc8eELLk0P/nTkQjAcJW2/jmD3E3qwHLnQmrae+f9IdAP6
Lz9ppcPJ3p2tf0TYFIx7qufuksFla8CNBKlNk7+QYIwR6uaZz1MTrYVOx0mEA6OCSPk8APuZ8a+r
xWRpDK37vK4Zq/6nXoZt7fmejJovpofd4Ogp5In1s8pQ7bcscc2rhTvE7Wzz1sPelbmBlBepRdJx
sa7b/V0d3J2E2K3jVQ+fnfxoesYwKTe6+L6Cwn36GOt88OJixcbC6+BQji2ajt86skGwMDYBZ1+N
ATDN1h9Oyp0ppxcIOfYvN7pyj+J9nKFzgrqz7bOOQlfuSTh7hdxPfDiQ1Z6B0FKMzAUqtKboNY23
XJdWq6/16omIvTEh1Dwi/AaienWPQBxVYguA1JQN/CwZVhEFRav6str287yFZn9evBftIeADzpzD
9vYL0gYn3Y/HNAJpbwS4QuknG92oPP00vTughc/aG3w7oYPfvNmLfCesJ0A7gj9uvOg+yBFGyUh5
efRVnZIsMKa/ePA9fRIoL1ENd1kTtwVjBs8afwA/W0mxLN27LTM/ZigCmbLvQA9XGYzsgN+Wue7x
3Qdya7nM56cz/j0i+p3xhEw5YHNWX7wRlHTuHfDXkWyZ0qsEsXh8CM2ZHYw7I/dLFsHG56rHzs2I
7IsnJhbwpgNusZolmZtzey6mUfG4HMoaofyOPulJER61hd3Wn5VsMkeXysypMBXn9Lj2v7d44ybw
QRUb58F92J1gCCOMO7ZDQn/ZtEmbVQpnGuWapom+nPKvXCHZJabwILo0skSeqeR3kbrsJJbTfUco
Huh3G7U4WZQCtCJdVDZTTnuKjw/fVqCbDQwB+vEh67PW2MBBXlPV+XI4lcv+/wVYowLRJaRljgd7
ysNcOD2mzPRWFwclXGZT59OATkgoQe7uEnGk5EtEYrHGuFR44XxbDTc/N84WVRK4PmZVSWEsw19T
y42oBZy2xAsh9+AHatvnw494N1OAFJnjfXSsewS/NWhYt7kDAplfxYxdbmrj7apLTKPhpkFbZzMH
gkaquPEaNND5CKt2jE72ywnHM2UuphOX8FFqWyDne4KGKg+dxYdq+qpzL0gDMGmczAa1AcA90kQi
YKAT89BumdUfQvZ0xat1R3PXddSqRhraQdBf/6IvPHWX+gkjkd7jbWbHUYzh+IpvcXXr2MjkCrwo
Ny3VnNsWUj2lqJWZCOYwyRr2XLWKwwp0/NRDJ1aPBhfUKXkx+Z9zJY59ckQpf0tC/qBqZfGAbqGi
cihdJDxJUfD5VudRmhEnHSIUbsduzkRtTF2jEEUu5ZpFnfUgQ8EozC2KkcR4Nw4m+1Nhq5pA/AV9
DAXWWw9HvWuiR8fl3iqzOrFPLk9YGhmeHCEHZJecNAPLiFweYucdj+2QwZ53+57DK8bKPNfuGjiY
/hzyZooOZ3NjiDe7NlsiG85rPGlBD1L9cBpcwXBm/f5XtMtihSjOCSntFNZnGHmci7BLe2FAq0wp
rTeUE3g3o+P8z8SEe6Xj4Y1/r4y2JCq4SoHwPMH1GBJDkdflytZ1I/ImOFxmmQTJLSEVJZnjN6H7
i8w8QAButErGMAL7u6g9382p/phF0kQDs3fqNPib86qsxO2kZBWrcHfUIEXlM56K/OSU+FP8AJzs
HGP0nBuipFdg09iVMhoKHbnSKlTXaotVM60A7IJAIcpNiSHrxJ+Lep9LEdWLSerXExZxbITv1CaW
3alwjReo5OS8tiKodqtrxXFfmjg0xxtb6n9Y3AfshoX6jqdPwokbb/rNK+PMGqMsXWEQApaHofur
jCtAtWG/BXEYjy4CN86v+gxtOyPvUS/9QTqJYObkL/Sp3fEsXD0yVPzbtQfbT5WB1P3pj+VB433o
OtYodwBrToDGVhJERWtVNVrwwo82Q9ohn70r2HY2xqTestZUJEG2sgFfk3wLUS8kEoeAhUsycVP+
tXZn0mc6q/9lByruscibLVDV/5+Z7lGa9DtEF463wOQHNidUmG2w7PQW+qtGYH8fVlGF5m/e88NI
HKnSQIOjLW6fePFqgKVtLyA+vY4SJ8co5hj6ASsy4quSQM9hBfbEZm77JtisTa6S0xhmFDtJkoKP
/c0V/2VquI/fFA+bPpn8sqi5hIsVfV1hON2bXl8qcg4rE9EeCkKrcn18EnN8M2WTaw8slG+Vlbi8
+KlNvIGirhWnvgfP7q4jzLtdbiZ+VPc3VairwlnAkaGiCHMUwbAYa13E45XK6TKtXTpgqdLxMIGE
+mR/Cbw9+gshtI5D7Mg+mwJ7snAMSH5la4AqRRbz6GRVVoeEq2EFDMIlrJqGAEiVfZkwro1n339m
p6cbm9ySBV69DhgbM/MECC8VfQDepKLHzdtExZOkJcXGYl/cu47CcGh9fpPkntDe9+zd7qvzHja2
Eis3fBkDUpJXIPWeJCZnakDSYvxeHGax5M10L79iGypSk654EzRlB5nbNSNQRVQckgKNg63xGfEV
lByaU/cB9wEXGLFQDWZHxXOUVXIb2JgQaKNxQVHDfGuaC3j+5OxbLRrvPcIXkQhn3RgoI0vWucoJ
eTmj58U3Ptl8w1G6/ZjC8GnzSX6DUVaMzbFo+YIDtZ2GTSeWRI8WocA35/Tbe1t2lexWNZ8gx1ux
EgssG+1sbFslblKlwhPjpk/Zrs5rzjyLEpotXx3Etv0MegaJ4KmAyetuJ9gDX1LkVifDkGw5idRM
PtOMrlXMc1zuNA0lrjTR6DrMRG9KMx4DGg/i3KviFBRa1zxl7RRJ9/5ZfwyT/hTQmsLmfTfgw+pQ
iJohqo7u31KMBUk1uFo9KdLnsc+5NiItSO/yXVuXdmFdHW/Q0IyG77xH0ZyjM7XCHajhkDOaRpsE
cQM9Zwboi7uQeRrCJtpCL706AXvMBBd+doASi+t4nEwtFBUZpSEpyPngwxJfRMm9EHjUKpxuGSSo
ygMT9jcuD/nwz2Oguacjg6zUeovYg0zqp/Hl5bCgYKPLIH9zwE3vmV8QB53arwaccrGE6tcHf/Rn
1E/51bOT43Vn/WLb4YJg837m7SDD5ikRh6IOnVZPAInHlBBxbLXL9JR6aibxvSN+GiMK1qZg68x6
Ud18KK3aCm2aLzrQLxg3F6YCZuA3udXtguHFxYK4tRmtZtbNgnTFRM+LkJRaQPZQ4Sst9YvpNcUX
jsl6frOdkYRkSlMTwBefO46JHb5NHpye/3dSqk7n/fP6JJfGYpGyZN9Eou3ZZ58MkNfgb3ZWRzVH
91broaKtx1zPkiqtz0sDwkpIv7P2KSOGm6JdUAWj65tCciETG/48xGtp6mK++z0sz6LJlIgBSoE8
JPRVaB82JArekN7A+wyg1Qzn7b9eiQEkGy8udS1lk8cUP+IXmJR9FruufqQ5Cgj8+lOLaoOelWGC
oWKDSh8zUW2sy8Gk4rMsZ3Nt3E7SwhHSy1QCVHCAPUsie2590ZFD/7h1oqJSLXne0qEKFwcFeFIs
MBqXb5rDCP2YjfwLucvH53dsBUgfYzqy0OKbUQck27nlXDXyRwFn9E5f1XcoYZ4kbj24FQKI8wj+
WTcODlmdwfVnk/ap49iEXOhe7YqR84LDd/WgB8dPqorZZ9qbSqfMd5z92/h7JSmFl9QEGxvt2T/y
1V4F2H7s4YkpvS0G20f7FC7Cls+v/hMSXwflTD06uzKITOEWiTwt+ZdCh8w+1V8ho2S8KepHAPHy
7V7TC50WmiCVj1VSCncRm8Ku5DrOuYTN3U/wxES6AF5dVFzKYDErkSySrjRgKty1NwK+AKGgTQEw
g9pQEPfL3xtCmdKo3sbCanxhX6lLh8T30IAzlt++Lez0gMejvDgORSjNIpqX7jc0+PgTrFAkxML4
CM2dmOP5yyCwI0WrbiRa2lLDXdRNa8/aarwIR3V6FDzIhrZH9Lbx/dB77d0PhGTOzTTQVXEXzeQU
IiGdNp9Dg6/LfrzlzAP/lglGKKxeMk4M+ioETb4S+I8ZUJEbpMd4ZH/8Ed3SqSJXDkLbA54wiB/k
DhmeJ7h9a/U2TafA3Tj5efNiZtzIGfZWzLTnyh+OQ3GEJGg67neQid4bzklZF1pUovcZw/VXmNEM
JjZGF1el6Oka0Nw3zdD8JlteSzLRMFyM6jiBjEbL8uCAeHavnp1yYEHSA297CjIqUa4uPp5EigQx
R4XsPIHWl9wUChFPzKRQKKA2oYdhSLSi4wyNZcnZDpkoLT/xNbGJiVkleztYR6t0AqpxJZCKnlZ0
zggUi6UXXok9pO/r7dr8lCXgZWwkOjRx03h0ZCJGIWCen/rSNjZEmAAxRf5wxEhOXykka+nvBZei
19xlVbRtd2+60j0zKsdiwLIcezVjihd1drRCopZapdVxzJuVRvu3TJAwEy1ScoZueVeGNJ/EnOrv
YMm3S24A+qwCyYBpWHHDAQtwgZRDojSp62wWMi1YMviFTiVHcj74BWSpcgPeJcrr2WXOoJhfdFeD
2ArxR3+Zb8nJe1LmO+7B+fF5gFrR9oOxNNMbRHoT58K/kHtWHvftWRL7Lpi2Z6agwT4UUszsmXiu
IOQfW5/fWVlSrHMJEj7KYthMvnSWgQK46R1m+qyd6uzn0+h3pej8FjovUE9JIr2YS/RR0r5lIQvh
1fe/29rxjdi8ohcgjR08QBTIKkp8K8ohwMDAHepC8PuFX5Hq+fpgrxasFFFUEMvnpLXm1YfHcR6/
dNITfYvE2PWVX/qoB9FmadtibPoaWMW0ot3ueRUV99EiGA3bkxiUVOhkWhZpCfE3TSLt3J+idCmF
B78QWq0N0+czAgjCK6Z+IdE1K5bXtrYskovS8cdma57CfGpCeOculLJojtPo1tvwVNV8hfA/muJ9
W/YkCUfXGYeyu0qOS4/blj7zFBITOl/PhFRjP4jQO3mTPVRbtQPQAxpqwMDcynRE4JWTZ0TJ1AeL
yh1+9aptazW7pBaKSVY2GDRsACixFLW69ZQ3Gz2ly/FbUJ4SxyrYUaSSAfMR/a+38LyzOP+e0QpN
WFYURe1G4FMeuHXC9N+6AB5kMs+ZpBfhmUF5ovhtaDhvKGKtzLkid7s99zNitJYYGoY6ws2WPnzK
NzYmMSCjuSfLxA5zZcFX0PeWgJSRdwfnY3yNyYeXOo6RKdBRWe6piBCFd7geM3RhQxfKOaN3wm7O
WYySy1xDAgCrZRJm7KkhGCU74q4YwbhSYZ6l6VOyNhGXDJT5sFyTTlhshu7QXSy0IRbHs5xeoiTk
H974nmhmMiBqL3iGK+VuEkIJoTEOwDvimR+n5dvG96YHTzlWKQCDNz2RNzb4TneRbcgl9mkDXvNp
fcQvinBdxlHAGxqyjmMrC7xx78o1b0Qlkux9KIjKmk2DlHeZ7gHncdZhp+Hbvh39zKNRrZ2Zi9HW
ylggGjS0WX+tkUehThvsuJ7IYBhy8y0cCKzhFmPyEVdjwyEl2SrP4PitLRa//W6V2kj/dxg8o9M9
SUwRLMZt8Nk8JCav90q0S9qGWMO2PjfdY6xkvZ71QfCzRmDZcSQl7rFZx54zncazjaeT3Q2aDDsE
b2KjkLqn8voBkdJnnFxYUd4dXjR1mmmmGrmNYXNrlfOS2yaebSyRVsDS/AidlShJG6i9B2xWUS3s
AZJzdfQSCq1CgswEs2EyKR2+uoQIZvsrguHWGXEeTGYBnRGS2vnD0W2oJ4WekdBd+oGj1wFt4ZPI
mcCZ+wyS52GB5nJx28uFVsFRKbRQJXOohTGJ78+dQu7A5fsq1IH8fe098FKW7Lj+olr2tOVJQDD9
7RKLR7kc5CqkO71FCAKB0JsUV6DrKAh9/eJEKwV1rHBCKV4SjqM7fI3ITIfKtnCMnYnNDlrzlHEC
IK1JrzbXtgT5nC6Ijt9MfAl2oZ/4fdi3cAcEiAUT1IxLwfjQ3if6KRKPlXyDLNYZ6UYSRz4UuyA0
+03zIJ3W+/DndsWCzKW+AMwDCjApo/RFJ7ncdytrgf7GByxtYTbLHF5CoaskbEQqMsg+Bb7sYvRR
qmF8NCvf5K8KF3tcBYBh3TRUrzsvkbtF1FdkXctcfe1nrKt2t2Ln8Lzt75K5HDe0nnT2qQ77kgcJ
0TOaMbQSar8KMxWDBIQzT9lGy605r++DE4RXESwQpQnX2aqikg3VwMeGfu+rKUXya8I841IBYqUG
tajbhF7wxYBOD6m/SuwdT92uNZgR5zkU6f9iEccRNkFQ4zJlopIdVq1RMCNR9QXkk5HwkRaO+Hsr
9VbuHorVmpZsDLaRwPzI5xFWUxrwMaK0Ga0HnD29bCTq3w7IqDGsOex/oc84Ho3LGSAkyhIbjsam
Rmu9RALcnHt+3b9rYem/XSvMGqDjVHNsDtLiYz1FMOzLN2ybWR6mly0w07mWyTmyJC2Q9KRsSMKW
CyU4y1mEWUL6tEMQ3qCePqL6pTjJNKEWj5PHUKP50oZ/NXVwBWCfth3jlpB4zXHd7osMToBkzDY2
7fQzYL8pItElP+Z6xYbWkcFAHXL6qhrjV0tLb1eqnWB8Mf7tKYrcT8d+YNJEd8Mqrfveoev7buXm
t1jhl75O2P4XKapZ4/HpAcAzp5JjgdcVtKkq6NSY4byTjVca8Vf4OhuqCml4Kbdk2+ukOv+7qGzQ
Bn1GXfFinA1YOELw7ddXGmfV4kFRchyvrZ584EG5/ENnmxKEFACWkKODU+FJuX+gMQrhGj/NkZXX
yb94NzNEFtcbVQo4XyxWntaQjWAT+mSjm7uNWYhDyofa/QCy8+GrRzzyxgjHTcQDBJGTvPw05epX
YNbWUh2mYFJWobYm4NngkeWO2jBo3BcH2pA6lImfCmO9Qn6O2BpYjWJ9amU9KMK1jtuI9s0mu636
QzsBCcv8242T7wkwathzmeZ2Pu/sOIIJYbSM43qMEQV1HdByNhTS/VEhLo2sE9owv5XC+T6/HhTm
yIQKkQq49s8EnB7EKzh3bxWxUD7A1sktFmMdyBc6HHm8dcuuoBJ7cPkVWE1LiARjioSab77Drz2W
wKRFby9bHfZRBEHiVmw71v8IaiyDKqoemo5ZzQgtZLhAR9np3tO9D6lPBUjIYTUKAR31khSM9XCq
fFyl3VGu0tah3l0rKm11vW6Bl5OLLFWAueoRQdjyK7a+u3LGLsfP/Xz1cEpC1Amlws7OdqAOM0Hu
Sm8rRIBZYzYEQkxNJhHA36nWX2hYvtlEOET03KFn+LLyZBEmw5ZFHrbcNaZprmo+Z/OXvLe4pVxi
tB56a3igQwbd895kXwnV+4wXDCAYJEQXz5DnSMcXneSVwxG5UXqfvQs8YowJj0k63RcdIc+CqJEu
F0Xv3iYadYMofia+UXTtD7HNzq1Yj6NzkeAivYq8FBy8F+8pFMP3deQdZ3Rrnon6p/A32oG8m0dr
V/eQNq+sW4+nOpHpUt5WYSR/KXDUgwO3ckeF/yG5dQGEWKnUHNgnIrz1/hXoIVz9xe90J9ImXx7+
F8KTpekYkyT6oXWKlbD432FlUJzu3VIf+uOIrwQSWDd2rQV8o9uCLE1ix1khrO54dVEZrgIlehVF
vN89K9Fr9PTPtAJ/Qyq63EdcJv8mU5C4f7huZpH7yyxnBKC4FQx57kFsyUPcCEp6zOmm+s2pak5c
2gpdpSFJfcz5kBDveuwW2kXmsSU73bHmt2GKyiC9rdKTbMbCIJ5o5d5RBR76V6ok6eJHEeRl3ZEt
L+Wab+TEU8XSNK+9EC4gimiStk11hHB+FyvzGA//h5Cms8ehFZbHazbhdwf+nWnGLffGScvWpCNm
8JwHSPKEyfsjhthLUD2TyFPZGPDXNQcXCqtfjhzDD+GhjeNyOMoPa8/rZFhDJsv9Kjsmg+ONiGoc
9d0mPj5AtViuXsmfmipR7/j5d+OsBaKz5IH/POY1x7iA1llFYtCJ8PxwqlIrkuteu47HJipmWqJg
QzrtIhfxLhp2CiotX3E6lICOGWfEgI1iDzWsjHg1i8wn7lD0xIqR5ZiWsrqL3LS83J/+G03/wVKE
5dCLlCbii07PZfqKkgxUuCyliIQ0FYUlq385yGOnJguDfu8NAfExpCfo7j00rEkAhg/MY+RfBSyI
unjyOK1AhTCUhg8gklAsEfnW6hG+t4zsIn9Iud/ixFurxu7w2S05l/Duym22Avj4HkKXlZogO/34
mvbOUcBPgcy/JqxXUeFowQWkzciqWkXNl2NJX0OWS08JSIgF3ctmIggMDVkb2EkfVkNWvnhUi9vs
oUYYFFy+/5fEr8/J+YM4hpnGH3dLOHak+dAcMrIKKiVLz71aH1uYRma2Y/e0m/hd96SidPivsX0f
UxR7hdOh0yf/F0TQVyPVYWiBLGPCMIbKGHsgDcoeX+COE8DXRi4/HcRxHCs1XsyfzbIwoZKHrTZC
iuYlHHSOlVfqW40BW0T7OrS7sJB/rYt8k2s4ZsUA3bQ9/PtJA7oL7+jFB8W3VLUg0xGj9ea0nNbP
LJ6kNz8UQ7XLwCqeGsLhSIWjArNsVYZGL4xJuvv72EVHT4ACqPCCcr3iJepX+PCEL2t64+HyM44m
Ewz2jsnq1KG+14EIpJchxe5TDUfR0dYZAof+mZt/tRMx5MMrnlr8/4YelLWVDMh996epFw1qlB5L
HyBjlfNOgQVYO5ID+UhjbTVJCt095+rZmoI9GxeMqSyxhTSmlfmvMh56A6Q+jx/Ds1skE+a0Z5yi
3wo0GSEsoqity1X1EkdKAruGNQMVgZB5U7ISzUDgcJapJf6Nmdpdn2qYd65B5lYRgkiDhrtytI1S
IQ0NB2u+CT8WuLjdZgl4krSDqjCxiDLO/xFWPT3g0fvkDgIaD7r4yPWBx25zxzc9M/icQMU5F6WU
gwhOcM/ShsCkUqPTYEB96SJ6fFbNXdKdL1pHK0s/0uX92VuigrcxWRPp4uzyewPb5VTBCKjuTnyz
911royJNmlEcWhSu0hSNm6QJQvgju0/EyCdgEyzKPh6scvy3Tz93V8fn/33i8DWkldidnd1kGf0H
HJJaJfhCW/rjYXiKJB6O20FxDE8JcyVE+VNpq/ngC9M6GpPbfb/k+LvbRmyGPo8p4kTKstcP7Fk2
EOyN07+EsiZVBFNsUNJxtfROpeoAcCGz06I3CgxKbO2GemnY2zEkxmzqG5A2cD/2bfQS3jhPVQ3J
zjEL1lt0x6fWDLW8xOPuyOlXSKJ2YOgTVU1k1cycf+3QpOY8yRQPyGssQOP0H29Ra0qzTDX2Zkbj
hfZv+AoDmeEhajEaPBYg76SFDHl+iCrzU+aDILyx/S9Ts1+SQ9mR7cQa/chvhLOBcP2KtrUVENik
HEB87JhtiTyJRAD/zbhjVlDotcUMgB9Ej3qpIXABgIUeNKF3zxikLxZh5GGMv+0CYokngx/bllwG
hq+Pv9a3ySv69Q3+Phlbvj05KcJYlY+8sJlNLonynywjG5YmVt5r5WWIrphbuSJyKOZkSMfacafS
6BLfZ68FVAYHSx3eBap0Pq+na0KGZO1cq9DUtzqvkJZairb6gho4IRoqf4GmZlG1BM1swmVRlVI2
woHTS6d67Nop+UVJ/7qcm7YwVW7MAaV1vHMR5A/4wm91DOaxBCkzXGGCkW+skBv3zBwUVu48fPzx
o1zcbNMVZxYLrENGxe2fBJPZlLFRq7g8ndvn7w/VJxRN8OlZVrKJjfRlGCiXDI8XUEBxbg6Apw6l
HXcIfbf6CMf7XYhxmVdIPayqyP5Q8B4E9pX/dW12NwFYYAXyrDM/tQqN2jwhI690Ej7DhR17R3sI
MyCIkIBzirM3CnJ3sxwShL7s4J2UtwhIEQzgTwfh2fmAa/OIvPwlHWfnVWRG92uQusCl1UC3mSa5
gEzxbTVAl2zVnT4l3h8z8MVyTKvHO2SadAm31KekDfr/6DEFFKVQ+z1O4YdAOyZl6SNkrqF2QeH1
Y570I8mFSHMyvzmBet6F5/bUFWFjLh9nZSML4/bUkn74JPqwiC7PtN4BL4x/P+E/hQpRhAKsL+vR
wrgvA17ngCovDA+Wccp4Bv4qRutYVCXMIUxyFrnTYjuMorBNzU6usw5GntABE8MGVnoyBn9VnA0A
/W2fdjZ3A80cqVjxzX59NNSGgW5dAkO1jSdpbad1saPctjZnFpMSpUSLp/xRJsYyA0mkecoshEYl
GkluHjLkz30JB8Oo+IJhEbpXVG6nnbnfkKVE2LfV95oAtXjOE6kgY3Grtk0uga4B/XE+OTXaNaT8
CB9F9xvLFLAbzoMuybhd3AzRLGFjODzY8WK81yRJ2KO3BeaVs3ips4tnppwxm1UVok6wAYn8VnSa
u3iuOVom0PGhYugXpoR0Lem9sKmvNN4fs8ZDjO+11wm8jMe2ZikHU/F1SNEc8lFJLJhcjPWFMvzX
9bSiJc6Ph3II+r5m33ZSlcjVfzai4inF2v2hlkSMLIot2IBW+WySctAf68SDOxtXbACHBjwbUYD9
Uslcehw58m90lQajjVY2TdBLYD7sK8vdERHlN/KnvOmmeq8yuLGgZhSaBRUlxuY/Pb0CiTHr4z+0
nuwFcIwd1aDZKMFmvF8sc7PAmJYGSeP2F78BQH3DiR05I0suCJgTTQ/Px1QC5NLVW+BkT4dphxWx
CzYU06vqyU2Y4of14+XEHuWhoFp0GiYpUqyENwnUdK4p90x61OEneBqnnby0cPB0dft0tHILkuTo
FDn9YhLG8isR5tpOZrIP9eciEoAGAdF05fabwKHS1TbQSRLCbRiSOVHx3mFfd6Vc2Go4/HswBwbq
GNYMWGhHgIw85kvCY3gvBDdoxg1SMlauj9ukRNQsuZmHqq3u7RJZNUQ3+VL//Fdb4XPW7kccv8Uj
b+DiiCnRl935rvMT4Q26kyulwxVikjK51kIDS28wOEPzYKlYC5hZ95R3vncL5Sn4cH3UtEc9HoJ4
ix1bYzBdIImftGVqkBsRBaZgceOda27n4zcc+cz0h9gntqAtuX0EvxZIQBXcLp0PPlVnPvjKOZoN
lDX86aDWpwejyQHAaGLd0AnVqt5zF0hq0onaZ0YNZeHcFT8MkqsIP/163Qz7RMUSHbIo6MRN3oCG
HqqHIuBcb9d62k6MRjw6pDko06iRNlY3vAoA0iXuKJUgx+5F+zID1ImpaClBZuD0SJjeldHkrDXn
kX1A78O8P0UTyceg9N4fDG1cmvAN07sKqT+YcPxF8k+DKARNNbrL0UloMmlGZpm5arKN5X0hQUos
yaDl1V7UykGPi/CLgHXKcNk//nSLJKj4L1CpiF8XV6kkNkTHaLVVbIE/E1Yv+6gMlv6itVVHdrlU
lXJpCLB9yRkfzp2CdO1TlbMeqzBaUUqL/XvVFTu0/naHnuL+KpddEuunYgChPoRliG2t8Di+Ui6A
gZXVTRlxgfihk99ja2wYpOFSMjmDRIO5LS1UhshP2Z2R8McI5Tru9RtQR0ROcMaL9NCbxKjeeXah
3olPYksjaYVGFKECx9PFOBRxpx4eaK/h6m1QilHb1qoaH5gwBALpiciutkM+8CgXbse0TgsExSsu
G76U/95Wxi+GakWha2fTCBTrWcXRaNOFAHh2jXHZkD4byAk9u4xy/y73UveiYxQqqjDsEydiegZl
ri9HiGzJJny3HMAW6tUZrOiBUX/K4QAWvSRvvlRsAIM8SE6Noz0fPVgm812qJTp0U70zfyL22JXa
ZfCIUaF+PNSbD+mei1JqGbITyXrhV1B/A3nYa3q2E67GRrakXNWc5UXASiWDc0k9MFaMwVOIvqee
LhewXX5ziVkT1IewODqmirAcaARdasId8O/TTRr+o5fWf4PFuxWawLqih2+RynYAMeHNENPMmjO2
83zoCQnnTun/Iyh+noQhcRgMsRD3I8EUq8UpsQ7tFm6vE7CB34JNM+rOGHoGYIikBSlRR3d3n+EU
XtA8lqaM/rgc1mrQugzuzUYadiFZYAgslqGcPg4oeNugXWO/UPUFdYEyOm1vl1at5/8vpN0vd1nA
cz0HyE/ucI+ZWBfZt/PwDdE5kL7p8zzmn6MCHTHCTv5kh1gMMah7LXltG/G1J5vg0RbSQOq2assD
G7oNMbcRDZS7l9iS9FI0MEm5dbeQe8hcVjWlMpU4mc5RyipxyOwp1TasgIaGGSbLMRNn4QrJi0dm
t5xekzqkJLe8DqJiecSSJm4YaZTJ0uFWMD53Y9siXKUpQfvLE8rkIEwWDiuzaMm8i8H5YyWKVT7t
t7dQ1xQ+zJlm5yBQ0ddXSW2fArOkowCIWhZ3b+cz39w8xB2KA6V8nErGLZODlQK/YfI9TuwodAPY
WWHjtjmidNf84TKNOpvzoUE4G/3wvKc6BwuS0qDLWMRp0YIjG+IdtShPxxlc5coajno0sf79Q+WW
XVIwCtLtKEIuvJdR77XbUz24NEwy8ktEzDPmmKzowsSLGydVYGNT+FqWvfcducUTn/k2yhhqAaZU
QO0JVo5z4T/jSEjI9PsmwlvHyygHwV7k1SqesWjvg3TjDcZu/PeKCmMwMLlzDI1bIjkLYrpOReDS
+GKT1+KWUpGdiWqJFdOgynCQ56eGGzxEaWVDqI4+f0EonIP+m91PdpPfPpiC2HYHYYqwr6ipFLIZ
kKyCAf206QxW2lfIqXt/uLrEc0Now2IXmyLmFydbozYLSpYL1GEdN8Zx5O4UK8aLoB6IKrwQ0UZd
nnfvNoGerzERINe+sXgzql31W0aId9iSpYtSy6v5BslKZRkrecHyOFWYp4BWxJCix/fs4qEuRBMF
Rwc4t5UivoKUyfU5bfLu7TpXaP/CWUVnOhVoD+IUhoWfjAzJyO2lvNF5whRvx+dOYBZI0KBvl0jg
OEsydxR+ME4KQlQuCunTdRZHCRM+E+9DQX3EqTxj6IY1OGl16rlyVLs/POEEZ8BAIiTGKATJMZlU
e9mBCrw5pOH0QiABboU3BJA+lkfhzzOu0ZokjQMJwK32xnbGSrU2zh6VCVe6lYOu5qETY8NNUo1Q
/MV0pv/c5dioLWlSVtKf3YJQs7+jW0PBUepbJEjr+Cw/edLQlkrI8TE8Xp7U0lKPVCy4ojREMdTL
dSFJcDfb9flIBLuOw0gcXMCuuOo1yku38zxlMlTMAg00X1/H9vOn9ZnF7vOIcxETCkFQ+4qktU+7
gbYV6PTR9wwXONzdYqkQ2XmLjXyYn+OvRBIV/grdKcvERAxENF2F4WoITrb+KNgnzNwvPdSn06hB
e6mVzrJaT7KEKob/k5qF+UDgJvunIr0o/S3g+XHRWP/BMWaDZPH2YhK4ttHNvqNAb3MXhOxgsEGy
f7otJceuVDiB64guQZCHdnY7/AQi8PoUjAc7ZvIbGQQrR0UJew6w9FzDSy/nQfEI8EfdfyJHnQF0
nNvBFNu1hyfh+J7+/VhNHOe/ixd9r0uJouQOUMX4K81D5lWsLi5As29uzBnxrCFIXSjPo6ScyIXJ
XigfVq59IpsvJne2c1gWmh6vzUaSHFnQuZ6ZAho9sXUNbEkDa+HCaXvlA7A2zSCWipZv8BEOg6XX
KC/Zzhm865RuhiXXUwjYMXoFeaj3zaou0p6+jh6XQgWJobGLALuHaNSW/QeKqRojhf3c3/nk5xLZ
Cam4d0XmKqZH08WLkZRuLh0d8hD+n6pgvwFw/7Y3gb+lITSRfCxpgx0AYbOzX27+qyoNg5aZwRpl
wMmG40nrzy/mK84JDbGrGIh+dLAdGzrOSZ5+ihAw/sg7FicODxiWGeP1xV+tZp0EeU3eg/DO85kB
wm40WWDsoLK0HeywSBgyCdrBMjlb+PGsZ2vhW782wbk2Tcfrbp4C3LjMLhEdDzaoD1SqcR9uVOCD
1VzrRHb5wPHf6k9FkGqn+CGXd6cLGO+DwuCDxgmu/ZZX0CRtSNiebAjFhrBdZ5NzF0AzliPezCGV
rIIZTxjmL0vYIp3TiYRPj/5B57roCSoEkoiFMEsBHjSyfWw6MBfX/5ASYGP8quM5aw3F9LDkXPTc
K6Enf0TYCJZdmJzt0RIVRqDiEIoNMbXwzvVYG15nkrXCOBFfrs9xLbMQ1agICI2XH1MPGyt0As5X
W9DNCjkGaaFkAM7+3iLQYSD3RnulAbfiwSU/DatXqe/aU0n3z2sfbp34vO+YjDgvKCYTAVNpM1+l
FIu0AOQyIv0C9exZXFGR6csgbrBoTWqwlOVX3aEOeMfoq+bTW4eH4r9hZHghNfAFypPnR23cf+/u
TW+kMpLWlndsDDDd2P2/8ZBlb6RQ+2mSvbSiTIRqENXaiSH8mMimPe/Y0b6Ytj/BeKTEUfWJQm5A
bkD0qIt62NnoTZdqkyMTo3N5t2I11nV+VtzIy5HVgC36oBKFAaoTn0qUv28lU+iVxZ+hj1kKC1RM
OR9rsV/150edCNGEGeONUkGr/pSZorl4nwsoKeFS46Iq64OtGvm+YMKZHSYC5bJUVFw+Z35gRR2b
bmyMmW5oh+/OC6purBFRSHqmOe9NAtAt3Ojmpe1aaQD5PeipEYyaLg8gRVfaPHggDYcYc0P4voMs
3oepHgkNNq+WVSdSjRkRbggOSmUZmw0OQpAtwohZy13zXN1M09oTTxwGo7GKYRK8DBtwouwPXFTs
tikE8c9ztShGhHFPrV8tLpIrLZkwtyQeeEmDwQmq+3s5qCtynsAHZ/NxvAP7xADHIjCP3AJ7OoGg
03m70+WDJ/EYZ/mbForCKNzeHH5p69pHN2wHbGVff8I/gc+6yephHaqsdpsnD72fTwc4XbRE/YfW
J8TKvhQM83AzmaPvDuaX6umfhELX3NBJ1M88af0GNVhH6SvyEUjoin9q3dH4pdpoKT9xweCaBlQx
YcwplUuurHNarQnsc4Z+1m34vZ1sVkM2t6X3iQTRbOaUCgjlD6MTLZm2q2FPRrEtWDn41nmx1iwV
CSIT3RJF6wQ7qkekI1MCYArvE4hAJpN6QxzsdktxH2qlMuuUO42tLQvno2j1DgAPfn0h/V6H6sPE
k8EF864C9FG8+H7cG6qOggCQGOSVQqUyMBtFEGbTluy1ZJDRZbKSnSrtZlsACw+D6FDprjvyuLjH
Y/cU87P2Smg99C92Df7j8y/GpssQaRGyGhzv1Y0H7FbpCxoabbJV9/WVQRiYzZL96iPxd+2CnQoo
ZVkUbxBXMXhtBgeCKWA5b5bsa6CafPLSobTnPEfSaTRgIANXNjIwYEuU/+FkO+PpkTJOOGHWecI8
yjhkTyF+x+Flwjgr75YEMJ5KKCUyVmVSODSaSJeLiXC5e6CCCTcSt+W73ngbscp4zdS+MUH1SQnt
VUc2Nw00/50ci248Snp1t5TLteow34PGK7xJMaag4T5U9GGcJUsvcgxJTAVpGVdRJFtGSksXHr/0
egTv2HTshMB8L/IZGgX0wkEXbl9DEZYFdeSHtnHbxuPodUnfExF1LhzcjOl0J3LgoPhUoPJXJdlp
PlLRNc+L2k6r0vBZy80PwkR4u8oJpJ2/08qI198DfcaRpP2srgtkcqCiTQJRf3KQpTDowTmeyeg1
xrYVuTJ7atC7/N/yubBrNqAq8bWU1tkrlGeSiJoQ8bolViBqAK2FntbFmgK5S2eu0uJq3EnuukdJ
kuPbWUT87JBoJ/VXJ/yFBe96bcwocYESz7uJrKQVdOVOBV0XLgL/U3UwedJjHUQKg3Iicm+/N5/e
PDTXau+u6itvTIygaAFYiSyAKctkE2BNbheXSGq6nqfK/3R5PU99X/sQxcGoExM29D2G21HmtmY/
qNay4vNp1U5D6B1GiOlV1vR9og1jJv2uxl+dNm8Fg1xPiQhFMsUi4ihG3PejaLGEGei9suvGvpYT
s+629uQzVz1UC9Y90Brec+44tS+LRpVEySI7lx/kFl5BLQPXTiJJEQr8S68YdmizaAq14hko5itd
KFMLqnZgCcYvsEpViC1gPZH9mFTh+ZsNG9ba5jVqKuVNHXD33dzBF3CojoWOVRdabJdvYH/6hoHy
a4rrKbDR9ol8JxAtowojAVz8GZhqlUhZ1D8vqfUMFlcvXdXbbF2EZ0JVSamjX/9+mZ+rzknRNmPc
OfwVQz+RRPIc4r7sRwgPUgKsjtdq9irYnXTj2a8ye4L8fJMDEoCcywW2Tcej8Vy1/8C7DPRqHJGT
tY/hWeDJOURH0B50skD7lCSmHCu9Q+QnhgH+U7r6VscfwfzoC8azDeZtb2rPAcjCWEDDzotZ2gIv
Fxr78acs3cRzC5gDW8t7TYsQT+17PxS00TDexCYMxC9xp2mGKhS5MR0Y1ECOv/7zAQ+fXdDZP3HY
RWxjiS670z8KqqCUlBjFLXNOhVG+hllWOYj85NXpl2B+lnNJsZ0CcgzoACOyUFYWGAe2usn1aKBl
m08MYptgb2ijBnqbb6jXe8Tnp30rpdI6FnhNv1KJRUWTQKUxYn3bPbaw+A/qXLDQCx4ySRF738gf
Rimx9ZxMerzliPdsPreKXfWPkefYc5xeUmRk1gQfT7ZMW71m6lGtEHQpcjrk64eYhyDF9NG9prdr
kPOrz/Bpp5gYa2vzlYuAqDf87zCq2nuekScqNr6NmekeK3XDehxzFqG49nfz82JHB2Km3oSWezsX
huOCyrb9m9eUSOkAltILdhksVA3XbBxjOKcC/Off5lPPJxU8K5xU21p6mPIJqdHmrzdq+M+8rGPx
N10FPA6ejdQ9pnxuXyPiATpwBGUeGFKBuyOo3T9Mw32rg4VxQceS6E2ngiKwzfu8RnXg2rMwLaho
GMTfGmEc1//k0vG4V+k5LgYPhwX0CabSFOmS4oPDU6ZiLIhjGYmwOKPZb088qgkANBVbgiLV0WHG
ASsh2ZC2+/dNjko9zadce9lLB8cTdobR2lrJ4G9ezaIzyZHoCIrkNKFohEJRmybXbMtKew53ZrHt
QA4r1fnY/m4oDo/PtggQt5Zc1p8N/BEh3+XPY4e12dAAv7mIVTkV0n56bdZ4y7Jbt3lPZfLeo3SY
G418tHWcVMPGid5Gk8wVyjJCxDTtYtjBIAPgooUYsyf+HZXCZZZ7Za5cGyhkvqzmgU5LaTjJRZiJ
Na/GCKS0+hH67nMh7TJm83IaeiJBf7U/oiyWKU+bStPlNY0GVhOa8YL/HxrKf8cOJq+ts4cE4AWB
iZItmW1PgXozDftvEGaXaeBgzPUrrk7Pnm1+8vv2cqXMqkTXfbnbXpep2BDEqSItrH1ClpVThvdt
gwlQ1Z/lx9D+IVWplKEvTEeSS/3Voa9uvnIW/0zaTVqC0qjpUNYMn+Bqh6y1MNydAJ0GEwf0Jgey
YudtpKK77N/Vw6lFvIUWpN2VrrEoTQWa6W9j/6OLUUKckIs68OtNuOYKR/je5kinWNMmibGO5yUr
TIWjF4KqAIzkgDqHl8Ecs/2MO+k2IgFNGPLfP4GNE3AIpUXtY5LRQDHlC27EJKdYm+34rwfvOwt8
ehq/LmahvKuRLZSZYIBpguf8or0/DmhRzhGtLphR5jJoiV7yyvrdzDH6xVtxKxftLji8eX9uo54X
yGZqo7T2pu6s6cCjMYNEdlgigwvbMUhnmTXDsPHTPD0B1G4fPSi55DICnwrCIJIGdF50lnG3PtET
ZCsy6F+U83y6DxpdzpX5qK276d/vagidMVLtwaQ3umYJSGiTYxMMZTPJgLb4EOJmBLxGfud5/cJ2
R4L3qK6jfcDcG4YRowAj3BmHiViwvMEfYDdaMLJDre0LiIudxsQmBL6QOeQkrXadm8ApuSgVMqCf
KWU62PbZuIPwQpAwmU9Kvz/jvNUSUH5Yz40Qz+xJVB1vS4BHyd2OvkMmNUtI7/uSfwEvuzc4TbMB
ykeKBFkimHMDRlwb0gqMxltUEU4+O1ESRj/bMIRzioHwH9pGIejwAdAOWl6mfl10d4QnMENnoR9B
xhMt2r72S2QqmciZocHWhVSYMB553rTgjgMmoBAHIb2vPBnP+fa06Xw0E10/DQyNeI7pL/m40BnW
eBFErpGVOyUJwHxXCORj2kXqir78byqg8R5N4UK/YVFRIFZR73Lv8r8SinV5g46/K1qgmyxumH8P
EkL1ETr4YYTves3zIjJAgAsBFLgLunjMcdGR1Dzw+zJYWLVgcxQPkYPNuyWRZIt6uGbNb6L1VjtX
Ovz3CIc7OeUnF/BHVM4RP1fcx64jS8o2HaWti3yE+0m4fQks0EDcVZtvCBhEOd7H06YLAnQ/EtY+
dnjzp4Rk58Pe209A5XraxyVzgLVESFBhJ5+0j7xZx26oaObvWtD2nzC1klp2k5CW9mXskoLYIOY5
6U14h2mDGQRJrqqlXGQHnfy013065caErVhM9EdVOy+PP5+PF6TtRow1EGBnJobUYxQs+iGl+ki+
H/zjHnkp2RZ/Oj+vhyfKJZvO0b7C3ux5JxnnkCxAYFc5rA/nD6CvZ4xqFXsq+o5aJ5Ko26IXVr2P
1AAvFzldGZhFFrWe/8T44uQCHoZpB4nUT8eqcX9UY6zca/aQPzPTy277wgIAF69Gk30vVj74pWVe
mlLxmb9aN518yd5CZ0aEVuu6KbrhcVmnAGYQrKo3vkpRTStIXaElnCOx2QoEs/g7wJougTFRQw3d
iY1No6FuZFnANjFPCHzmxJ9tgt07P5RmtykjkiIPJhvastuYJiK8OpyQqSmghFNtUA9s9EKT0z6G
VI/PG+EXyOM4C7NQDvY4d/7DG0JTaMNBv3xurI/FU/E7LNe99io9OAv3/aUTOMDpk7Sdg+RkI7uI
RJruKkVFQAACbhkuh3Av7WhgNHWId2243mM7v0DlQy4hHHH13rbDN71g2aj1C/f+tzUC9ObOfp4w
YzitEoqJs4NVhZ4BxZf/KeeV+GdDxuP69EYne+zkRYrEw24NGp21vRVAJzkrF66w5U9qy6kBoPTd
6rlkbU3UTdTRpNtwjQCd8MEXdbB6Yju+IIHT0vPEHOEg71hu81COrcOiJDXlhJakRxoUza59Xjjx
5mX4JEsJlxAyIuQIn+TY0SYZ0yWAyLKFjGpUOkWx7c9mngCiCK81ExwZaTwRf41W1+i0vsBDhuTo
svAsCFBQskqt+l87X5HBL9i0/SeirCQqmbdMa40n8pvxsxrn+zjyHmzZ095IVwkGFvcbzhHec/fL
Ja6+WzdJCYgZE6599h5uqMg9aXjJ2vFen4IoUFTYK3UYj4WSW6/hHtVfGXqq7ByNPoSoJb0sTZ/u
p28FIrB9vG9Av0rutOF1aYQmWlx6Ao5LexJ54JCuwGB5ahnZSS2eDZ9RWy6Fa9iNb9SjgXNDVvMn
StrRse2kasAcGDsDDRt+Y+HRdUnWI+wv4t67L3lDJc3Q+1pr0t3tAwDriV79hjakj0J9ZtPhDLpx
+R4UJC1GEOVmxdsm+NWOuOlb1fdIo0x2rJHP1jwQ+o7aO6JQKrgaQkvUKTMd84Uc28ViNqlvIjyS
rk6j1Jet2ELO/XQ30Wg3kOgmwZrYCoOz64vZ2+mWV/A8XWMie9SX5hnfRk3rAk+fSZf8xeRjQf3H
HpoEm5gJny0hhcvR4Z/v/dzwO+30lFrSLc8NFmKXSzV53DcLc9JchcXDOlDAUxDT4g/1YeCU0NCF
ULWMTvrLCYDvql+xYEGJeuiOihjAVtZVPNRDXsfIBVbn76DiAU/pwCj/ouhMaVHgXJUiJQVwa178
xtqAdwovGHATSAWnbklTwKMtCw6XtCUvTtxjB9S1ZtdNyCHA7txfQb7YhlEA4dvw1N/7fmJPZlAR
1rOeWj8j06mTI51NmV86pA0IUWoRuIFOd7sLzMY0LoyVqYX+aVbsIco9J1dHunuuvO12Y/izZQl5
Jv94upL6C0JNG49qT42EV5FSzuKOdRF73ouZpDTr64JUmBHcXsNwXw+rV0lypMumJGsG3Ye9ILZ7
USmq1bfDpYYiuErftRyVdiIByibtAr5f1HbD3g+GNgJ0Zakhc2eHZbK+IIzdmZgpaQ2mPYtJB3xP
lrnJrmIVeoPyFErrQ+iJ1FNJWt+JwUc1yH+CW4lBkrmNkZVVjMtneWEcEFgjBI7KNkxBywc5MTXQ
SszpwG2nqiun4Us+9be6nB4m9kULSjlMcrQEmt8SbVZJgVQ9gPe8f9JDPyWmdp+0vhJurMnUN+vP
/Dzb4DozNF2DUf94k0MZR70EnmH3Q7ww9OBSjKE3v476wu3UPlvc+Ran12FXrqwKxK3KmJjlkZAE
LcVmuKoCvpghCYH26pE3r1rBk+bdJBfrroXlRw4XHhXpiBL/5tcSNtxt/deVlITjvLlLfLxYP5L7
u0mOHMhHEjrOMGFL9qESS8AVc/thA+LdGXPIDVSjp8+t5ZXvKmEE0pJDLWEmncSiT3+mB4GuBnMh
3fhu+Npz3ABtXSP+0MYZBamjH/qw+wfMVrPf+aRo7qUw8eguJ3s6QMLMZ51wQA8fb0ji88qw82Wd
DT7FZ8FZCkhTozxKs7wW/Q/4MOxHgPZkMNcRsyGOnR8D9arCJ1BTG5186btXs+XiI2oozK9oHOcx
B0agsuM1MDVOFUGAUoXmX4NeWJmWYxqt+LJwbU+L/nRBXZUyde22GfvLcNANvizzqnXFomuwZ+TI
Yn3vyJKJZi0FQTjrJ4ZRgVlLpQXxPE0Pliup1lJndBkDpi57RYO1UHrRRBGL+F/BpNzW7k5EVhm9
867/DYSqc3liX+QWRzgwijd37XWeHmrDw9xKMLMQKnzniWr0AYPU3N8rTtUghglddei91c87yGyx
+VjKLek5pPOEIeM24lX6Jw814mJ8Cwd5Bi9WgbEY1taDjysNeuQyfT4PzRdncz+IEabYNavRPMbx
N7nNQGW8Crq0LDPxof1zGZtVKzp+wOmTMh7v7r1fDRqyhnd+23iMyH5/pc1851cT/gdDSoesfWE6
Y1e/qHCoiTlG4OnOIb9KIyHnDwuVm7qlMfsLt/Dx57bM2vrehy418ZyIy9K88STGU8g0EZEjtFfQ
MeNc7xuhf3FBF9q2sOC9ZyOofTDYZRDdnA91qZTrE4yBnV3VypmE+5I77oIlQkF11qLaAC6BSZxr
zY1PpEDD6ip8ygTXD29AU4xFdAWMYe+ClN/39Fs2t5NNjDjRcMncRGqpMTs2bZ4hEw5RMVNVjdpC
PcJzhRgqmo7OwjhdWF/xPTBGRkBovvVkEdZt53Lg+AgtS4EOWJlHU7irGtE+yEVYRbivAkuh8rOD
W5azhE9DtqhySE97pI9jE+srlO7H4FqFyEPJcBHGupf/3cys14YKrLlijIm+sCz/93BrdZSynvfw
m9SiuCiwc9FkowLqNGeHPnL1m4XNv3dOzWExuDJHiEQAjv5anMVpva51rnK5+s7bJXfOYUGxB80Y
XJRRnzCvIOwcUkkrMc8bWwXWTwahaZ5mVZTc1BJuwvwj3dXxMyjyF+PpvtwnkL/mRV+ufJh/rlmU
hzXKltxxUDs29U+FrEuke1f9UIiaWSav8lUXs8BXJZqXqti9rgGviV3qwJ7zZBZB6y46NdD+nsSw
R+FXyr2gAOZ/4MCDbbAwX07ldwFR+bRFcU2/kOje1PnU2fHyPKZZ8pUPZjozHh+5hbcNeNTXJqvJ
3odLwoHaXavJZFc8yFYAB0z8PvOUqTy4kodDldeyclXfEXl1sElXiIIdhpNYf9+yi2u1TQu+p0cN
sA18wxB0v+v8eZwPWRebG/MU12rWdIBJs979ZeTv/4TnCGaZBaRR+ts3OycMRVoR/SMTCaN8fqjJ
7wqK82+w733ZR9pgeg7zkhgHefyTavR//N+2zMxFdfbNRtyf4ASU9v6zSCMvjSZg4QEOmnVZXujb
iuSnMWRo+GtFVIpHHdqcqwluyFGeiB9BFf6dIpkQzj8DOKX5o1H9FWhWnQ+wvUz5jT6FCLh/UYPP
R6i11Opm9HwA6skMz30g6ArxYwC1wDWQiZ2pfjW+M6QlojVClQjHW+jutsbNS6TCQv1DARNZoPnP
8ReXg4kutZxeGVbw583S1+XyQ+59Kz8GLwtHd7NHf30EEfd8Fho2rGldwRPai+oMaRErg54RPoRH
j+irPOlBrDePeKZsUX/IxbE/AXques6bsqGQIIt5sU4Qdzxdb85myoqpS7bgV+LAoQQQrZnhuMY5
hPfWJfPjoWlPf20tgr6DIlcS4SV6ELPMwTMfImA9hLJMDpc2A5JLzRyct2mnyzBSrmef3qSIBVAK
7OZipwixna7/xicRkPMsFDnk84ST5cu6Y9BYP0jUTp0HDn9AUA159+Yy3oJfCWKfc2yHX9ufNm9p
U+is89eHqrqpNJS9g+d7I66+WE/VHuc6qJN38YscA2wkC2QyT7psmMiAfN4mfGX0XVc82n8tHgtG
A/p3d3UInvXVw1pgQsFWWc2PioUUfP/+yKpJ7aQsK+35WpoBJwjOGyXA0c+D6Lf7YEc2DfO+Jpe/
3nfACrIlZTOf6sQio7sFUMbLGlis0be9T8xEevE6R1NJwB3Hc6pqp7cg4ZRt7YOHG4izh404fl/M
UGM17yXJFQushn4X03l9dmVN9XyxfRl+3o05xl8X8v3k+yDCaxTy/FVM96gAjKaKZu3fl0raVGHO
fG3b3eQh2r8eS0WZUeq3OtC+asRyI39RSTFVOQBlkWF9jnCO5jcCxptR5EvBHiCAVZ6pmPeFBBMQ
LytTz1UYH7dsUFcKOGehbiLpSoBxVjFmdAL1sLg5/xB22UhzKsMQYAWsMmL7h0F3gVQsL1IOZu0M
UnC2tdFvsKHkRiVSmb5/g/4Y6qBrI7pZR2cTbCi+Sb0v5FeNdDCTdZYMPgEFa0cBENcTVso3JdF3
jRkFauXD+OHeScOyAiHUB8wrgz5Ad4YVsyvWiiL1SlgO43hq7CVva80sY5Rgcp5n+ZObuYgnsTuq
+PWcsB+WPKNVC8u28fx8bAMMNbMojfLXfhl5iME33ZMa4casQ8+NBA/Owt5NBk4K09pCBoZCUCQx
Kk6mDQIyOMxTuMdIu825FCgNOdJnS7oTAJoochuwW3A+7PaFpFcVXvmi+b0slTMErkUu6xQ9lfjU
eteJbZPNUlmcL6fXFRCTGJ8ZZCFL5E5Ee9Zu/uHZWG7NOR1+1XCEYVOowHs3vaWrQr2XqL9rSUMA
gl0tlvRfVYOcYl+rvHTk1l9CYpRl/PI4TF0v4idZZK3CdkRJ3N5JBF/vBs8GGIJEQhQAMWAgZAmE
s5zXSknbuznQTUDlzg9bN+sxvGWAxXn/10GTPswcXJtnwkPj6PEltjaBKkA/7+f/v1YLN3MhXCaC
gz5zyK1u8ZUPfyWQ88fB5aZPsUX4wSaKQH3vkhaOMClio559vwrLkAHNInJAaBxjHyfN8svU/CC0
L4Go18IzCg4FfZt7QdON9FCrqEKyCiZDmWqcVGx0ae2yAKoFDqW3sFMISKuC2ExYCa2AL8jTt7iV
M1FCMaqQqqjBPmWVl5HQUzWraVnScdCANJbxQBLkcFQZFZNzqOCJFE+9bReMjKpazi1Y7Rt9tlYR
DH0wqDOyvutVfAZO5Kfb34ZCOqW3zkWd9FpXw7Kc1nHPHu64M+44x8o2846YVU7bcKq5X2iGjZ6G
DgzcA4f4VlqIolmMObNH2F4dBZ0dJ+WzrMrbHSHm8PBUC9l31/+h1wV5/8eNgPudy3NJyODAH0s7
nJnZzwfs8rwmwPXqsi4wGzf40JPwQOvU6R7gm8k45NcTMgNdFEPLRD3qcU8pqktruX07xAY+GQAs
o71yJnJTpNu5GIFQHqiP/L1WTqqx7qbMBjcYv7KNTbLwko8qHRU569+RApm3xG/MlyRtJQPnwoa+
U4uV4XDsW3A2KTU4MbSHm1aQby8J7RxXtCVOcUPfey0ozXjbuTvH39OYq0eWJ8rbwD1kZ+dHBoUE
jKkXAi9gbBg4J+ugnWQ61S2MTW2ZDQMVOruPICI8dW4xdwF+V5G1Ek1iWCMthP6xi9Zh8SsKIB/q
gEQDfaCe8T0L5RiVtCkY+anYkPyW/BkOCA2e9CuK429Kh3cVpLuPm8gFMYogholvdw6N6H9c8iF+
Zxp6Nhk5e2vC7km0TvfcvHCyR5uK9Q0utZfEMDSbPD1Gzkkg3RfsX9RUzyo/PZODEQekAiOp+tJ8
Re000/I39C+2EoLJtYRW4R0k40VfYP/RL3oaLQc2XCcf1HUTAKiAKoiNgrRrfZYYoLqPcKmkCFBr
QGr4eWixF1MVmBpb0MvwehRGGFtWt0KNS0uDdYnjjLDauxuDcv8RN+yJqTK7cAomBKoKtQ+p7AgV
BPDS42rffndQsHwwQCCmLFcqgYusY2kFgkxtIHK5MhBHAfp9YQtdx0n3G9a3Rdl16Vbi8ZCmJ+X2
NOZtwFmemJ5E+cMr4m2yWJ2Y4/fqecr2+8LVaq3FIoKEAEJEy2tYaIEB/2BjAlJpgSS+xj6UsXi7
SeJlj+i5hnwlKVvi6J55g0w/jsd+U8sv8ppknh4MCnGUak0xf6VmIfbgWdinaNR5SwEEla99ylzZ
3+HYP9k6wnnfEt5RWk5ZnQ/M4Ht8X3PPMfe11ewqKLOBSNXz0ZRAHBVlPHyf+i/HjXeVbrYPYNsz
SEIvKABck9PwnRvUAOQ+jOu+RAZsVikoCvn4e8PZQGjMU7qGrBp2LatVLwfnwimZPGoSoGCsCnGX
c09m35r9xbGd3gcUfGJyzhLy4pMfReKcKZKp2QzNZwz6NATj27vNKvC/n/kS+56l65MuB/J76qAA
QX5qD68rx1kx5yOS4kr8Uv/QbqkPXul5PGQH/MWtX6IMvJFTOqKrGryitkQax8z6aRokjlWPX8gB
zAA29O386yRiD75moG6MDWIE6Nd9apzogFkysl31ccS1/UwM0yQyCjNEY+NxSLcXGG7jRBXfNw7e
13f6Yu4mXG4MZqKxlQ2JSYQYVN8kD59mD97rSDj1Twg9Lrh5Qp8Wxg3Iisqw+BeTMh0wHPnJD1e1
AeVj4GqgfYZGOYqZkcKSA6liW4ZI4S+Zv2LeVzFL2Yk3bBIrgEvr2P1U1UwyNjdNXmojSU9TkfDA
ltUiFjGPE0rmaHxh1KRTIVCK69CQoo5O3pCdA/F0apJcU0CDhlPPkz5C6PWueGlykyTJzJLfL83A
6N3GK170uOD8bIadsOkiCWiTBCMCvr1pXHED1TXN3TGI4tMbFFsoY21g1HSy4AnCH6NlpaPxXb/3
Kgnw7R1A1LF9wKv4rr2hEGUAxjqpERx7dgs8ATEvog05QN6i9P0oE+l7BwZWfa3/PGBGAOqTWHMq
arCg53YRLc/QtofBWQTW6vqcOIlT47FxwEbC25WKHXRwLRUboRopbaySCDQmElD21ECg3Guk/bKv
J7kIR6lwq9oj2ztb1CoSrprBYlVvYA6mcjBco1hdmWExcHLygZjRcnOfT7qbaFkweuDq27JmW7bx
aK940d9g0Hb9PtEPbwMW6ZQsAMAqlvI2tMfRTqGLCoqJktoAGFlOREnU+xWD2qzxxYDDWVERWppT
syVemL4SJmoYIb6a+W2MlrrFQMML0rrlr5iiFZNwFvX9vhPdDpVJRLuYaJ1AMMxLsTRAWWkitRcq
//RsZEucmhDb3Y9obhc1APns1tI2DdJ+AQYrYYXnXjf9JomWk3Grp5HpEbeVZMvhgdcoauc6cxyd
+aY9Ch9UzZu7/oqHcAXUc2RUldyho8+aDCKzWS+Ra5LXRcIJ0j3IVJldXImnAKb411mn61eFyOk/
RV5u9f+65wacz3SYF47ZZdoVxBtJW3Aww/qN96w4m0dARNHOvwfAxEL/Fsnml5dvQX3ZywEULTCE
1qOpVUAH5R3wOeVShrWYns7L8y4v7CQm6WaHxhMXBs9yoHiP+liSWmwS8kok5lJDRf070Raqr7Y7
EiKtdnFEgSpMEYOirzO3cZqoLqKUco4Dfo+8pj+FMs3Ag/yWZjbko7GLYXRZ4M3Y2kbp/IuyUsoi
u45DLY23oC3lI+k3Z31j49AEdSLeeu7xeppHU1HXVUlwFyxAzd9AAwIrN1dVj1GgB18BjX+M9j4X
eJT+y9jvEfK/o8esUAAIuFi7nh8UVQnXZyrhq5mkQ4sce6yNvkBEqfA634Ih8GtnQol2K58sovZt
HSR0/jjB+10vAH5zWyNJ3IcxzyNfTWEYzFF7InAaN92GD6u9hEGHsw1p0dZkpMvO/2/aVB8XPIb4
yfxyLx5wTM6iAzeCUbIxnHD3AZei+rW4hpSbAp4BrMM70cnnlq154I7YAiO0rXeYIJdhivXod/Dg
C00wipIWmCSjyswbMhLGSJmxm5h+bzQ2n1WIXp8iA8pIlKXT54fAYOO292Zzpv6uBAkVkn4tNIB8
P8LNNjE7LXiNws1TMr/7BA4ugurjWFHU5ShjF6VIG27sPmaKCzHwX7cVpXZlTKmM7xYhZ6+xMrMz
8UkkgXnLZQsBbiKEBLj3TwKNzOcryPNraOpg758za0cqDXGq3rot5pPdlTVvt5x4PYO/8AveSXRY
jDbJlrEhEvIigrxcXDCNtYd9iRCM0C+hs5jjwTF3F6Ts+ZIdofyijEugB3t4vxT3JxebqZF8uADS
6Zh/kiiUwWAbMiflxm2xTduFVR099TkFFJdUGuqf0SzC+xq5LzTxdm7T4yg9jGXhQvhAsAu7MGuI
M8hGesb4j+Lp4WroNROhCtyn5aNGrZHVvP/OqdIbww4d2+itmOOYNoBRYs0m2Vdk81+jYTFI1jt9
I3PfsrzTt3wV4AkBtDnb/T3Wu6TiIwTheLixijC9ZXxvPG5LXGxAyB9iHopcedo4QuctT1bc5OAF
DspAzPuvDjWfiYMdxW4OzEbN6pf8lQqIMfqar/Mad2aU4IbHlJ+vSw1LZOInC6GGoLafq+i4cUo2
z0Rlx5i9FW0ZXhqKcWlxM8Y/Dw6nK9T8Lzea/ff6jhto2v8gvx2LVTvw8H2aHfMX67ITEk8FaoT5
5PzFTQ3h0uuVIq8ZvWGhtaTw2XeyDZDKqUOPs019E6HiJawQ76gFa87PAvCzx9M0iO7R+dLJwZzQ
1w8ZfkTn+3RaSYcQb7q+soBZmmCuH7rV/pfFb8ac0NacGwKOth4XhhIg89HwJEkA3azGZpn2bRxV
oRNQ/uGIMTKuO3pcsrx+bIrNPX269SskGLrQNt8q2lN1NH1US5etA3Y4I30tCJifJtX2U8n9qijj
tTA8Zv0T2XfZNUOne13UlZGFvrMdkpaxvfoqxOTbNrkOHezwE7xb72Wib8z6kS2vl7fX6ZCCbL7d
zaXoY1lWY5g7m4V538ujhUeughuTwkFbRXrFOpCW1UTXQWKUKQkAxrSNr+O5b9PLh9gdb9Tw7TIW
fOdlWSpgfyE/ad015PqafCySNp+Dk5IrAyU3kGi9SoKsaBvDgWs6DNG4ZAHp+i5rJovvk5DgzYIq
LWxckNIEJ6bjUOJsguL5gIs1a2qBYfcSY7NMi5Sb8xl0kh8DFz9PW+HJ3IL4in6THoMDT8ZSKHzw
7XOKAcI4gv+/AXRFRbc/+AJKtDpm6/WZ/KAi/CPC4N15DjDjarGSMJzKf+vI6hvIZEXCV3doXFvW
dLiOuM5T2Vh03WSWgrhTSWOQ47J1WS+snBFQTRVlo8g4+etJYghrE2V+8jz3XTF+H/s0tdQC/2pZ
uNsqgyrEze0HR5+9Qp6YGGR7gtMlrJAamCWJBIyByb1JAXV85VUgsfAgGScl2BVOztLbHWj9q+uA
VUTfQtUw76E2y91WbjJQ+uifmWEdwd2u/gwx+juD7C1jXgSscWdpDIlVJBHEb6qYx+U+EJB10Mu4
Snc6NLdSulwFcTZcMsnq8++xp69fR5P23vG9aplkiWIVvXyU9FFjgujag625KDfuevxKE0Unz3v3
xOURugB7r5za7J5BwpVnJC93y4O77iUTCTf4Wdt3URkhrskG2Is31x3U7ujPcitqIUJ6OGqeF/sM
2rSKjFq7KK3K9P4CtakEILsBRWiLs567PacPf5a/xWUYRmco3ASs8Eo2l6iq8R65kIj6pUx7n8PO
aJlWNu0zrXPKnhvI4UwMbgEj3cqVeS4pkUC7S3AzCy16uG/3oS/NCR2G4T8FGQLpGA6i+E6SqVCB
cPpfZvEPSdQz6KxgHlkl5PDuO3sFGn9H6fHH9cMXXhtxNQYtLx9DZKyUKnE3Tod5EUY20oj3wjTr
zLXN6qf9TJlZmQTZ9/FaksXAur77fCKvzaRb2qLAi17hzlhiw7Lhxw9xQHA0j2r9PZBat26JjxOy
JbjnWdfmF8jav3M3gwocgkFaM6Cvg3sCjGU6Eb5pldGkdvvlcZr8C1K990SyZq8XL0IoJEouiTk6
VrPhITlBNByremzBTU52WebPGjCd81C16HOx4LM/98WkaXQHSllTKlTLwmjbardiUA8qh9kPHjOd
1Ie/6wYn9bMGJIsqs6V4bt5XaaZD78khigkl/5t6+4z4R7RBARCfoDtgxnlnz8UrgfuhHNB1LXNf
Zwu/rTnR1O5dGTF0aRoFdHK23K9n8yUjQzzdpC0StFQiSbZsDEuH2JW9yYoPVZTBsSuYhWM9XpsF
LFaABpOxwEWf1aOYfs995aLgM7NcmJFE4W+HKUb4KKRb3DBhDlseIrpPD1yJ8oo2Ar/OKzlai8qE
cGENNXigAOsrZtGvIzN2Vu3Fne4zB+GdGhxThcInHPpasiVX2IY0YUp+hZhAW4avCRgkBVbnjbF0
TFbwTW0mHjaNbWDNya+cravpwmEipgNexTw2Y8bSN3JhY3fS/4F3Jm6vUKS0SYofbGXgYwcgFMbP
ruyatgbyU2FIybiCT0dlK0E/YDzpMg9dnXHWyDjrs9ILRzBP2xkIQ6swdfrX5Bv6BOtczhnri2vF
NFrYR6WzTompFTCZgKxK0MUfx+z0B7THYBcvYRTw2uZtjvJ21cua3q0tdomomZLZyyEZk03T+T3v
b4JVDnNjJGenB86CC7GRIp5iZppu1jDfOjWMiqvzcCpSE96d1+p7OOHJXMMTXLqYUCtPF2cSY018
NIX/Z9KT4Esr0q6VqsYY4pn18ZUt9n9aLJ2fuU7cjyoQPWk7a/NqGIzrCLGY+JqfqCkppNZN2wGC
wmDsWNMiq7C0sRHr9Jn65tA/2VB1efv8WS6sNCcKvhGhbnxxo7YMhOjqtts9xIvYgqvCTgoj3DEE
ft7Uck5AUJiOwMraBsQnLA6x5BC0I36fiGPjY/p2CmZzifwghiTsnqzpRjnKJAYUoMJS5RdGhRsK
8y5NY3B3Xso26fxWvPF36vgZW8ou+fHZF15RZqojFP5zYly8yRDn0IuDlqwLDPtknunVXCX1vgTW
bJHQRyb+Ox++RdtjL5FJ7uBCL0x93PvFE+DPgSPHslFjPuak14QxELmngBkO3Q6McyO67PGbacXE
S6xHASfdr4+QFMCXGqfXrEifbKYH1a30M5/4Bb492FLPdo3TAjhdO6a98dIiAUoE2QpQ0UQoprEx
iAXxs6woyGi/+FiLor9xTyUCOMhMjdti3vTIjxhaUx1Xv9YTxQQq+NKTeMueW5rtHfx+VkWAq+0U
hrt9CtOWy4vwVrH0HDQgAYQRo7cqfkLjwHcmVGhfaG/f6ErbNLp+nPzN7ek0zm7VW1jXzMM1egij
qkXVBkgkLZPdrCYV16SG/iofoSHQ2AE8JjaatZ34th3xGKuTCwfl5++r3Br+41NcGHoAiH5wCTgM
uo0wTDrXTInXeVYn5RosX1IBAdvzeBRdnjGH1kWYjCE1vmRBd3RAVr6SHkWg6C9Bc9t6Swa6r3Rb
ZD6ph8TzKNGK5fkPlKWwyKlB15gupEAw5jQ83AmhgX4FzcV+GfXNXQU4Z7qstktg+lJddo6rIv1c
h8BreND5i1CEAGlxxenc/nNgFYlKZGxa1aLg0FXvF0NTKRXY9Aj3bixXMSrMqPp18JcoUrLMm0D1
o1cyz4+3g5DqTg4uwfSeZXjRS+uShjOA5fFRFU+0Fb9XfWG5EpiDCM5uWUYJt7Ev490uvRGguvpp
mBFtv946xXd2eXvUANAlPB+/wRw/n7dciwBetk4EhR7bTMwUQ8ORBcy4SdC52M6MppCcXrVnIKVi
iAlPLip+HhrRPGbuv5LOaYXMMQqDnhj/Q/ItWzwSvpN29fDcQWfDn4/GExEURGGcQhtBGCsMkElF
sBeRmAWuX/URGCXvc5AP8ppAam4sOuisuQmpSKS2bBzhLVVUlnrL/NH7BfcX68HzDOnISQTxQcQE
paUGkuUldmOySRHVVCEE/DMJtluSxPDLudDqdCQJclrDfuWuU9hcWB/AedzDQMz8GTuiGEOcT2/z
ZGAMxGt+Bw2a32VLGU4W+5fdpdx6YUB6lNEHmv5cxM1PBr4Ou3eMSmxmJl0jsg7mZpRN1BoQOFuk
M2rAs8I/a1dshsnsjz/K1da0ofBQlZwMUURnJAmHoEzsK2wYoFdLFWzkWGLltM5grGfyjSYaE+vu
3JdicDRPAw/cLwpr15Ayt77G/k0Iztz62QdrgXMESfm357iYIwoACuLJQykKGgvKSezhzoJ/06pK
FMHywEnUxH0qOv3LgZ58a9iqoHSIlqXk7bLR1CDtNEnXN0W584JiXaetZzly6hQwcyBIVFZGWHb4
sEXPGEfhXyKuy+bfKIHS//ARtSw6D0YWsI45Cngy0xZ5OKau8JBrvOgeac2CwzYy6kAoNkq9VeFi
5e6HSjnDV1AEC//itvGHBg9M4s5dlR7l8CGwGGfaW8uSt/Aq7jvqhL6fkLXm/xRDqYfTgFPeAFYv
YuGm5xqN5CAu5K42gXwdMnrvIU0pfvDxJb6NphTAcGKgqRoQ/JFtJrlm9VCX+WyaSMvONC2opk3P
L7IPjtzdvwrmclN4xDWZnhjH/T166Z4xqMfdCr/POgm6/g3lTVIJdoRpMX/b0j0IssY6FvnrRU9B
ig3T42l8h0oXEgf1ReU4msxQSWFj4Rz8NVGt2sI6E7JFvLMJUhE0F5yZcSt2TWPfkNhSMG9WkUe7
u0VvPbGxplKmgGWP0nK00I7Nv0zp7Mtz1KIPxHLew3AMEkQU64VT2nwsZKmNykNYMrNA5QqWqTSe
BMSRQstDE5ZvdrHt/6NBGSU9feFKQI6VHlDTgmTFlgFtDXoioXzIAQ8Dt1w9k+LNkWcY0XQfyX5Y
f/OuuZA8BDFvaVvDIvPK7H8h1gWDPPvJRBM8yAVtxjgx+oZsJIPrWVLmbWnLjSQR4ecYwwT7pbQ7
+/5X+ZZVOnoY+QXQX0d5T1PC4Aoh/wp2QEs6FT0CttHTa02wevI03g2/7Ycq9w1rV0Kvn15jElth
SaZ7bEOT1z7ivKhmKLwXG8Ud+NPCO8okfRV3HD55e3QIiSsptmKF+OSnIXS24sLuxzUZS0gpf49v
UMAXCJX+8U6caHF4OGvf2Nwmweoj854YPDoIZ8nvWR+h4xNbbQC2WnyoVpzPvOsMo8ohQAmWRYEK
0/64PJC1Elo5BSyUSAGV250SAkOJdfvJs7ad9sRtZS3/VU9S73iqIkDxEDjE3tWOGb6yoSnBWslP
2ugxS0I45YZHlMOgIl3JkU/L4q5x/l9tP9nygbRoNZFf9C7FwA3mMa/6Re/zsbA6zFiqjCI2akpf
CxjhscwXROrHbx4uspKc4+lzFn46u7LZmFiiJOD3o6KyNX/iy7O17KV2o8Es/dV9tH2uS3xmvTYY
EWPk1Ic5ThGi+WfYWR6C8o+jU7KLRSHX174VdiF1bgPMx2A0R/Tw8VZ4WTcQx5uUAv4xupwfF0oJ
khnl6pL1ObfWAbv6qxhegdlaxfQ6TWqtUA6/HewvqETxCFaDR+sH/1uXYM5QgMkc4FyaNjUWVlqa
wlf1ot5LVnoimb57AUELRLwS3ppRSL2Dsd2TkeOMWGh0HdcCgVC/4gJY6YX6TzghdHKcHZIuDesD
Hc2UXhfM9UcKNCaFJ0yUgEgkXMW5EOu4hh77k8giZOn07LAic6KwzBWEHetcwTreQ3fTDFt/RSvD
mxViHB2PVZEHR+mIlqGj4TVMBuvV0Cuy31TwRl36wWHg1qBzT1i7DxQE3LFJsMExaiCZuFbBhKQu
TySQpwPozDtXTWHD6tPqzmTwkOCpr8z4qaSZlnFZ6n4vPEeLKLxgk0oTx9fA9iZdGbUeKntrIk5Q
7ujYCzmvPEnSE23vtTg+S0AvqRiUu21vZRRwDja3BUgxt9wRezTo//w9V9OOsjwNu9VEan5BVZHv
hbibhHwo8ezppo78lPGNXUcv/wd9lVk8V4ol/YcS0ZYVG+MSLvCfC9P+dHtrHV86dsWNK1PScIGD
Ky0TtJXuTUtRX4GV61e+YpPp+vKxrU+AhgIno/mjcsxtkWjgpLgXH4D/6JUWSzqmieZkWI71y62g
NboDDzfdpH4PCXZBL0W9iSsK2FkPTgBOCY/OewPDGVv4Vp7wo1VRl1R+vi1vDXM+ayJ5qznngayV
XmLeRjMV+J/TnC1tJOD1bIX9NgPth3/SsUzEbRxw87emf4yfp4GOE+tda7XH+Ew/y7f3twCbsDDZ
ZQz5usEkRU5HvoUNT6/vTuVcAoOJ/UFpnmeD3EOCnJbYzKDSxdvEK+wVc9HjC77UzmHEOHoXz3A0
OMlU1IcDO5EXDH8jHtsEvSKp0h0y8FvZsw0a5upn9L4MEQ85ALiD922lpl1c9ERxmx6T0k7ZTF95
ipjKsB3Xy2GMx+2q61QdaVeAEcHI8i3ylQMyfX1NFWsunlmTgtJzvQx/q0oO49jIFrQDHc5B/eko
yqVsmoRmyNI4LKOBn3YdLNwEL5r5hfHZL+wvqNmdsaxJJM4GXjWBZ9CkcGqh0RYSdmrYDH41Jb0S
RA6xvd4wyP0SmuKQMYW2wlvNZXyxa+o+ypZYIEB4EGUNuHb7djWX5lEqXQ/2VUsEGSXD4Ajahhej
e5hJeTsOjmDg1MRj9B37wylNVLMjEAOBoG0Kb7gLvYXk8zeBkaYuqktutyOgnDq9cm3xRKvPvTaQ
f/0LbsgqXXaCaHkm+LTWpzTIyqztMmjPdiSn4d3qdSNFZDCUkvOvoBkHcvGuchBQQM4/mdwBZ5jZ
xYPIWt+Tr8Qzkc+8LvVBtjUlRFhdfoZzk3a1LgrtKeHxG32vVxPv9RHH3JyIn2rnxCiOldD3IfTk
/G45oNqUp1vevtCY2d8+UDMhyI344WvyZBmuD+anus2XEhflvhS7NiXkHXPszfxMojKsiXY9ex5O
OOkdlyyXPbKovgIgj2ea6Wpc9ByBMTZT5aCh/wzuwi9swTCj+SBNLu2o3BPIKntNZuZQswpT2kb/
mRmQJhV8ukHzUjzsOZqGmukGxJ/CiwcWEu8VH9trUvVd97nGTnYrZx5TwmTFmCI3k93RTKa7xmBp
eiODaMdTmvjgNWPWE2pt2ERr5dLkoi0Za1Aec9EfB5ri53/0lWpDFZsVyLXscO+aqGl4g6uuhgJ6
NFsDM6X5CUE5tsy5rQkLnBWr1aQgV3b9O2T9lHqFdq7zHUXIEpSkUoaNg39L4/bEuhVQ5PydpGVB
semfV6EA+O/HrDA0RABoOOkkDIFtCVZ64xR4UilFexy82fvKiw00+KZzU1QRHagYgiAjS0gtWi68
T3tAZC//bRkDTVQ1rgLz32TZhHWFTS27U2bU65RQNyWk9pSpgwH5j/pTNeTLJcsXjuCCs+ZlI1bA
0ksS1e0SRbTFRFclpEyYwElp6VJsbnh7jDG0x6D+qXYM2fn7twaZDWTHczcejClGvOwzm309dPci
oZy9SMvP9kgl0PlyQRjIO8e8EXllQsbRnhDEQm+s9FSDA61WE1Um3Qg4sgFJcxZ33uGzC8OpOJ8d
8fY5YdBPHcsoiKnFTs2PcD++Qdg9MEcx7hOAkJj52Fef9tMS321+AB1yaZP3O/BsU3rfc8e9xZjf
LyaPnLjBBO/uguTchTl1RoA0SQS8OeS75V/P6xJePfvz4LCECUxa8MQAQsYFM6OoZaRXjatPXzA2
Yg8229Hr3M+lrYq6p0zCGUzYKnXAhriRrS6lX6Jq7Q60yTVibXK7duAo8D/gTPLWwcJ1I7T7bwZ/
+MS5Kfe2IC7MYshhm4YL4OAh4NTIZ3NECuF+k6dKHeUvz3+JFuSgIYPqY1vkHrETYi84aH1RCbnP
1yAqMNaVwas9rqM/1cZoIoj9eMgDMGWpabWlCPnE51Um/fPhDbG4C1AR5gBHdWHMbsp8b8+kUdoz
Ldbyu1/Svb8CcC7QQYd9iWD1yJH/Y8AndlIHYuA+k9Ce5azImwJfsCqSpwo1brAteL7URENP1bk1
Tq/g+OTh7j7TPAjLj1D3lKZDzNO11WVjXHT/p1RmFyRqGuNJAO3uIsyPD010fWUuheaFNaAe4x35
mSgYzMGcIfjMfT+qFd9M3j8i7X8J8/F83QipgVbGiqg9tuGv6AEk+G5w+vD3JoJkBrMFPIrt6nLL
RXEHE+44Kc3ZAO9oAc6dbytBCVrz4hPleVw1HE+ubxkggfGWJWKXYMbMN9X6GGEt8qZ5jsyJuH72
awgzRiDFgqguh8bm7TdWCkpVvSg62Ebj5pNPt+uvOCCBovIJJJphg/jfP2LXm3+KJ3vg8IRLe0he
+Q6oM89G8loyicdfIaj7UObAbK7cSf1BcgAB3bEea+rPYrPBAHWScXQp/5SMINEnC0hGzekYDyrP
seF1CwSu5SolRFMuhnG3fhGhTC3XkgxMuNfgXFRK/Iq/5WOGAjhDkJXJbwjwxtfbX8v+l/eKcZCp
riazj5mpXhGucriZfxgHoQYVx0RleRN8M0VlKDlqywaHHwK/3t6lunvNyEt4LNHBgR+FlE4qsB+n
h2Bw1eBiE/mc7C3PqSvwHSUqtNpZcoKDKZQPbG4IxVt8jC9pfuxgJXDDsDwGw4hFvP7VYTofgrXl
44C/hf02rPPRdEBDqLnOGlOw/C2F2O/KuWtaJLsPv9UfT30JW4UBvVCN8dEpgedaCjjFcIvBfUZM
6GLksbdtiVqamTFlNPBJXj4tjWZ6wFglH3IxW0oQzs7050TB0YxGyTht8+okBqoKJNrPh9Yxvbsf
NTuMOe5S3oRQkvz66e6uOYwdM6+Y0WJ/ZjiAVZoWZviIyj9Wj8WRmkj5sBl8WV+gY76gNuImAtCs
uxsMNR9VaY8E72D9XuYvNPxPaogi0TI9tzTA6suMhLjjFnpy4SNhP0UggKbnqQ+h5Gq1sYVYiD3y
Kgfi1oLjXf1WPqZBYVLuDZbCniU4RzjNbavJmAnw1TGf+Lm2Zqk0r++AxDZvlaNqLBGN/rjzG7lW
RSlVGq0QaYVndMcrvUBwn6WbaI/ikXRtSQpi77rmjif+trlPjUP/ZVDn82AaEOQjdLxIQ17t9Hv2
jjWI7TV1t1lH7EwvNU0vzwA6pNIsZBFnbKUWCxoW8TBT+h/Q0LOrwO5l3v16qgkxh4kzkhXpRC1z
Ttog86c1TX0ObzskxZFPnltzvURmg3tNJZqjdslylbOB8L9Fls+1fcFmo/jnGOzqY/DNtdg3k9HL
6Ici0kRigEGLiRDaGjDKIIdLWk8bZmxVqR92wHD+UG715lPJjGvDr3kYS4yXMEdvPTw+CYkALiw3
pDhUQSIXaxWVmYCtxGe+Je/yxfFC9LlhZ5Q5mReJ6mat5ZUDD7uOmT9gxOarOX8I28UfXTmlsfv1
Gr7EFsF5/jEKArDs/Rw30702hYZO1vM7e0ixK1PDxNwFX2+N053nZmDVYbX6/TvmQO4s1FR8N1/E
dwtbDMwBMhmbHceg/k9mw2MTVqbxFW0Lwlg/jcwYkFL84cmUWm8UILDrBxGLkr3iwl1Q/LZvSRih
lYoru4eVZGGhgUnwVECsOF0mS/3+PfHdhO/U5xgdpoIC21eCPJaaF5XD3zPe3mY3orE/ZcQRrKa3
J+l9bECc6lrUkGIX1sSCJEn2iUkM3MfqUuEleC1fLfGyJN+ZZK4yFm+hnDh5JvDoQPZdWPhLdtjo
oPNnOta3FrMIktTZHFiEwUG85yYpHv3C52Fb8wzBxrMtZsC0AHvIS0BIQZdOB3c2+egBEyjfkPIB
oY/AIOmq56jQfP/LO3Z1KGxX1uGXXQsNFq1kn0bNuF9Mqv2OJznH9GyRPOsadr+7vOjRJD/dwdZT
G5DtLeYIs7rLH5zdMemF2XBxvID56fNZS3+DmnyRcSeF1Caycv8S+JJDXq94pA1MsGVABujfZgM9
jQL2L4Ss2Yx7juhgtKV5Ihp7CNGX09lU8GPakK9K8w7ElvhvFRv4n6qLoj3mJwWBwcHVROKW7bp0
yTtRA0wGlP91zwgyacfudFaEpIFYcnxyD7sB31Sez3dSerfkxh40CClxmIjpikBEuZoFDK2B/CZ3
9KKWWY+Rd29eFYnpQI4uizTbd5GUNkqCsfoWD7fXGlbh+/vNrpHH5R+DjNVDRugSbPMAEbnF3zsg
M18V9Z3FqvyeC71qHPnNWM8nHzfZRo2mpPZ7g+LATR8vhPnGJRlIau0e9Rqn7B9ukAZPWTo2OOTQ
oVPaMlRG8QFxJATx5DIE/gyGV243nd8MRMfF8AjfPwVvgNHfukDo05IRT+xNu07jBgLbZjZz9K7v
XbyKEJWJKwHLI+1tvsJna26dVGZodsdtMhjW9lt9CB8mT/8+qL5V5f55YuVkSRJq5Djo+DUUT76C
8R68+fd+fTtAShl4YQdv7+1BQb0XKmUAtqt7eErS8VAncFO8Y5x5o1lX/wopXn65kcEXZkDNRt5I
AddN9HrecmYILOXYtxuMi4qRrpN7244RE4pY2rym1jf+qtW/MEt6tYqpsFmndSIjKGs4SOv76bp2
TqJcoTTifc0G5WOGKC+XEMGJe0cv7QZGW6+UNJ9eG0d+PXr1+h2rg4ojSym+yrJWIL7R63aejnOd
ibs44klZN8t58CKfzkNw5tcLPwLnJirWG2eytj2HvkR76+XI7Oy+Z52Nokxr6wgQyygK7STHmWxs
+PgpgdAoNzN5B0pdl9vtd46393g9ZfeOIZD3Opp4FbkamAxhzGAVOOg4Q1WA3eplRGeydcS2jWTp
EVdE2O6HJx171x9qsNIX2FxDdRuDAkpCHoAQr75p/9KDFxUfXnRaw9ASFTb7Kr8Kaidb2dKF9Oaz
aKUaKvwXhO5q5qu2/FcXPNNNYp0eobssz/4iBUI6xsDQjC1g+hKf35PsSgx39KDlqAlGhy0uhcxX
gJkuuAuQhIw6On24J/VJD+B5mPw532lTw/MGmG/5+OVnRrKEvaW6ekOKdTPVoGdHJgW4hHIv5UHz
92pu/0bkC4c+zTEDU+VL6SDx9fSFcrHNlsPwHt/PqAsJ587DxVAy4Qthe5y8H2I318uIu+daauyA
5WfnI93bqUx62mdXEMvTIbmRm49SndGED4KQG059mCkgdwDG6M2lRZ7g/ehzDDfPvG3lQq8ESrwN
k1qMy31LlBWEZYqmm5ORuQxtWl5IBDGXsasqJsw4rHTVfj/s/+iqE7SZw/RF++n+9jjiqloiCKt/
odBv0iJgJOLR0yYLNUC8kxufCzjoEv11B7pB3atorB0rQLmYL/inIaYCqb+r93wjaewNB/aa5DL3
w4LKky6n8t8zrLVi+sIWiysKtfaq5Wl8RRlYYA7xUVU440DllPN1iuiPiLLu3hKqbeAInwuYzPLh
cq27sGsMEuH9LtlFW1NxBV1VrGemfTaKJPmJLRcIfQme7ashB9w+f+h+IfM1052MkPr9chuJe019
Hc2eNzIcuXS8I2EimeXJlUkLy3zHPexc9UdbAJnO5VsBi3Tq9KcNscLx7jN14JTM3JVzIacYNZCz
uuaglTsx2ZAbI0ABpfZDVqiOMbKphxnKXwBHOi2L+GpqkLoOEwT5hV8F8e1Kx0exNytRPE8iLVkV
gaQepRkvEc05X6WAfsGQQbLbqd2VYf9yoHM3M1lYmnPqh7veDSn2oUblJ6xzGrW3+aSPkZN9OyQY
T4jEa0ElkozOgODA4Kdw9jptQBGlosHyCBLFIthniX4tZb/SeqGYkELCMwmP+9Pu4IRbL3zAVz0I
dt7HYkbAFDJ5EsvAYfaDWVuhDzF/MOhNovIO4U7O8sZaPXg65qaIB/zx3DHucTegk6HeM8dfpZf/
mC7gPUYOu/Shwu6pRZN/kUkfW5NqbZi5oCu6CS7iXmnoZsXPTO1VUx0ysVax7thA5UZYsYdnzBWs
5myLFT1YexCXnPPGBCkoaxh8kBpxhwNSogFPFWTMxKnq0oaF4Fc/uCJ+hxZIa32UuOPV/vVROup6
z+ns3ELTV+RRqnzTlcdUt1VU+LE0TMVG//cotObuwjMZhCu2SjgwfG1ti+gd2GZOqyetlIsbWNKL
fntM7zsTbrwjD13homQh7zp4jHSj5q3Iv+VJw596HUK/RIosT/hBGoiwYZplyTv0DSgmhV30/xXG
PPM/JgDMR+Y2xTjWtKy+ESSITpHYXjiBVCN0M8rcM7WMDDHjp7ItN2LO8DS/90AiRTQTzQ/LzaCS
Pt0MusRBtUy6TpqzLPe1ImmUvUXVtpiLQgJr5uWECTl43nLxCqAauW7lPzibwkov3LbDaSNMI5QW
Iw5lGowrfrCQAHjdpCJKB76tjKMU7wiJhsxdKldgdtXICAduF+TmDZ+xTJeUqTB6FTAtuT/TDztT
2nFqUmcCkWNtqoMXlmPvmc09f6QGNUTEIEbnbffx4uj9wEVx7AA1nJUC4n3wKoD1c/gJSy+VDH3Q
rvUJozNpIeOEFWem0OFcvBrVJRXFYyWmOy3s9KLYnewLlKDVRcSdbR4PuHsFB3p3bcdcAv07KelY
WrfXaIliZxya3DrOQSvyWfL2V0hh6CyJVwRvhJ1IeXdLKLWuQz+Xj0s/UiymTXi6UTiw1YJHslLf
B0qyUAcVwjozWVymf5sVzVC4aS4WTSJq87aaVmIEGbvZxOrVqEFFjX6aXYbX4fdg3baXveXVSp25
U+OcADEIbRhpiS0fnXyWC34o8HS7KQQUkgRQ8gI1Vjs8U9G3iw4fu/3pHFDDdRFpScHnc/4iqPPA
+vWcn/o2gtnZVeIAlzdGrh0G7+2hyKSDucRp+2n5JTjT1cYrV4DNh7ykZIiMAt3aa0BRDxwNu8Xz
D5S4Ns4WYI5E802DUstz6X0WxrsLHVA6koPIvDUk+WH8TAd0r6499VtAt4zTwE/BeVGAZtn2aHpX
69rMdnMNf9cKQwzMbfCzdk05GsoMrRQrpXmeLGw6Dotf0XdW2DXS6Xibz7b+Brair0v5m1LOZP1C
G27P8YUI+Jzq8xgJwb4BhHy6E46u/vBm+tK3oo04tZjXB9OMN+fUzN5gWbHAg9F7q05N/rdVKAIR
hNZD+B7NogI0HtGqqkYfOk/Fn6eR8yjYIkM6+s6diB7ALAbo85NCTiaUPDVXjqaQjKiGF/bTArlQ
FmcrQAVPn/KMiDO9QOhhhtLLLb200437w37MYfQp5eg/xUp/CzyTYIwBxq9Zkx9/G1pLf1ul9icP
OIWRVOegy8T6duV2T3qoI6wRpswklZiG3sA4Q2WtVoRjNONx10Ae/preL2gRI2BZARBIm3gWbqYO
7o5bKmpq1QM75HVVgHVLoROM/fpAlbqsKsX9yJ+ipQoMFc1gmiassfLeLVv3scEYxDCMimwFwJP8
TPJGWc/To/FaAUVktck+3gsJ147ZWpKlmpxXTpGGqNnNQUFG8N5MubTiW1wbmdubTNgrV0HsEUMV
N/b9EgT/fPxTaW76NirC1r572gPl7rlO5sg+LViIuojKZ3zidLdXDg7MimDhd5ne0n1SWHISPvlP
ZAznJCx91QKy1Auy9duF+bcROYtkPdN2FNwAWNIC+PPSNhSrAUrgX4vgoGEJhC5G64Ip7F435Ydq
S4FwCETecbAN1avyvTLr0J2MqyN8UNavk94LjBN54Xw8mt+wPeTos2/w60+towDwaWJ8n6ediz+A
i3Dzc3czIkenCVExsoWACmx12Xzanq2TI+0YZwbBfIN3BQSiFnEM9FCsVjMqLoR7iC9IbZEf8976
xt/6LAV94VpIuiuY3XOVLlLKUdsvBifCZV1SwNvoJ6fzuOXRlfW3f/e19M5EsMrNTFWTu6YYtob7
BREgL+qgbLmeuis4o8R+bhOLJnjvkuhuE5nhc6fGiH/Qg+fIMxgpcXnKMDP00H1W+SvJ3KtuIiIT
JR2CrSQk+SAEczrljJCx/QUSWY5AH/688HVhIwYNv5dntEZo4aLuEv6rTRBAIcgsyHZLhrk+h5YB
HxF01pwDaPkfzCNpU018W+GhC67vkA+uRS2WEGHafErFuIf+coHYCObAi14GumMTFzXuq2vs52QF
8ZEb0vL6Ifge0RgT6fFYlIFQHClC2sP/Af3w+W9JQCxK/0AoJv/XFPBlQwa3wOObAGCfSs2QFD8v
536SVak40c+/76y1JAyaQ5wmsIZivZHv81JZo5NHJ6pN9RWHk/iSIVeu0RFMhLgnj43Cp+4EtwXb
FBZHb6mT1k6vcTrTmI9/4T8hHK2krhQ2045SwIrS5GzqOkIOzqBWA6HhFqxrpETknIaMOyz3rGZL
Rqnm/VuDHwqQFwDPCmgaSCb6mTiy2dB/Bsx6ZqxDwXEJCd/jjpxOZfK5xlOGZgCVVzJmrAx7XA/p
GVitVLZEkQeqa/zMyTv/oBO4t11MVGmNwlGt51lV/fj+L/LUMo+9YhNnDuUzXW+WU7dGlFTavqUY
jzBnr/lTidkwLwJjMIjuT8ljp+2dTrPtEb6KN4OZLlsOeGyk7E7Ce0McK1etYoYhM//uGkCTIkN6
bYo/rnqPZIt8MH9FWcbtcyubka5218ubRCoMRqg9gUX4SeNKfcEaqiwf1ZCdL2Me7CBJgjbaf5Wc
V4trrKo3RKHK4mGQe0t8iwXAhSUQB8gTcRc2WiLq9cMI1S3KgieviMkjZr9kR6/BkARyatCeTFxo
0l1+ieOibawusPxqaZVQB2i9sKIrU2qkiXLE07TFRI91vCg0UYUcxZXpNRzAzNdeqTW6Fp3A38Zl
/XIkv+jiUPttD+llXVb/jq+Q+W0yg4wQmA5jX4RU0OInsLD3Gq0bEZRVVOu9HWhQVL6gGnc//Vtn
9dStx4I3C33TiBcjTwMSDcovcs55hVDSltdHHYZrti3SA3NdgIkk9R0Oi8iU9cEZtrwhD9+BuMRr
P9eSoj92UDIrR0yQFQ+KjBLHYfu064hRfO3UX6RNgIaTuVjkuzCyMw9ipV0zFue9yhOHQ5Xr+D4V
CRijR+5Ro9yEOFhX6BZeKXUz2JGBlxTsmy7X4mFXVrmRIMANh2BIvf2xqLdrkgBjAKwOC3JMMxoi
5PEKR/2yK9rJVJes3hn5N+OGrEG7yypgNQMoU8VPoik7nQFDHw92QnMYXhSvVhvr8ETZ1njqKxDo
349f+YyQ9oQrEpUbVYkWuL9yJblPycb0MF2hNAZXO6wNP57k4hoTymiqXuVZvSEub3mnbPH+4+hi
KbfAG0wUhX8LndFi6Hp23V0dm+q1FYbDvwujCjqxP2m7B0QS7RnkT6O9T6PfMT9THifnYvRasf8G
bf/lnnk1K4XNkrQTaya89ci2tcGk2E/oLRHB4OpxPGyu1eBG2WFiexEUw0Gya151zMWlARSOki6W
p27e4wwPiTcQkmvNmnitxUiwwhIgE8IpE7IX3eA0+kYZ59lLcRW8J9b5uxLB8jNziL3IFz+If6RX
Gh0SiPEVPCIeKZj7BmQfynzUl5ks5HFfFMB8PLvS5sIOZ81D8tLn94vI1hLkBvGMtuijGlE+uzPP
N7nZJBz6FNXquetInfitnoaP1yICnl2wsQ9H8nf35qk8oq5p0wluiRdCGL1FQvuQPtRauK20Qz00
XSNxXBB/0KRjBlww3jvg/xmm+Qkfgd+JUpVNhcXcVLdJ6bjr8LQUFFUGG9bTzxbpEQ988kr4aF+b
cibBqjZfrezqPRSQaWK5HD6+mWsbfz8ko3HPny7OqA2W6hi8f6NIF80sO1j0j6nCmgCGsZaLRjRl
G9DURNaPbQd1AGjo8kYXBIIVh8LcUwx+bAp0VOYbubdUmpYRGPKUr6BgHvMISgb2ETlum0lXBS2f
PbppS27Y/0JBNWALTbo8hJKJTLDO8WvVd9a2ZS2HeBZJFhxKMoECciweBe1aW5+GHh8ZU5xJYAZT
r3cfVQbWGCidJ3IaPNZBaCa0Z9CffvejGoAGonZWAu/1Fmz43aj/T6s9GsxBPcL4CdY5KQDKtKW6
PKL+YHrwhCsyzlqlx1hmv/zhul8zhsl0A6nMiGxv2wIxdgvheNXEei4RIQOtCIhnmNk89sRlXuGf
aQB3+QHlx8ZZ2DjLcOCQ75ntcM8oE9kD+g9UDAIAw/YPZjE2yNqzTOwppdb29eBvJUleMk4YkyqG
/rADhGOfB4ssO1vgOcFHMG0T0KQxnvpYMhmybaVCKj6TVVpzk2tvlDGkTPz1FTD9cpzhXLPfjUvl
coPJiyU1zmtMqO8SEAN2OrdYL++7bl2ffdd+38Ng88gCx9IUc6Kyv6NiIKYZ9t5QfJ/qhMT8Uh22
24oWMwUPVUmgdNRjCn9Eqw0CLdzmGQbQYd/kP/8XaCGoEdwH6ArYpFqUT7EKfWnO/T3XIq5XbyVI
uOpyIvSRJq16oIjMxOgTIUueph2Tkcr456RgCLnRdrfaaK6dIws1K7os+czCvCPgFKVdECDwpvAo
mTNrmf2EFleUaAVXmkLrfUdyaQ+sT4zkDbbE9kGj2aVAKTbfpq4QHvnIcwhGJEDwHgmsS1rlKFZm
V5vvU5lNmo6hsn6/04ECQF5SDzO7CXzwszaUdNDongtdXcQORsRmd8q0tgYnl/OiJpD93QrMrszC
Bx/9hNtzheIlMoNr+tYtYLxjfNZyC/hfzM5kAR2O86wmggqJkpzKaf1V7+HD/na/LVbmKGduEv8b
ujxRewfXg6cgYayxWtHsYKkK3/DcJZ/W60SDrnuh9PBxRfIIYabMHOijaco3pQZHp6R479A/5oil
cWAsYjk7uVZk8q8bxVxp+ek5Gr6suoZOUSeYWnqoFVvGlATG0ZnL8ML3Uu53UEvqeSHBhVYkf7yA
NJijKcSwzG/5mpOi0bHhptb5vNeeikHt9dhAHIV/qMqkfpsRYYDlcO8UURB4ZAdhqiONE3/6TBPr
ZwzQxXacr3ubvhLS72uiT3FiIiOhEgQjPLrAWcpChzVZWLowNosNAZR4KrtQ44WNX4kQFFvZYMWU
Eh+nSKWLyvSWDtwuEZgvByFcIFbzMz/5HrqiiyN53l5xWD91m7oe50YoZ4ODTs0IsHcei1Ajrem6
dYq1ptQunFDw/c+MjzUVBgcEyuXKZ44p506Wb8SIKXYZJ0+zXoiWpeGdLmIJl8XFwNVnbtuUJCng
1HKvrm1IghEwUCj3ftExLszUeBv1mLYJjT6cHpcRHy8rDeWrwYqh2sXAiKI0s44oRVW1pesw4y/N
TBlUyTf8Y2CDfdHK8QKkY5ah3l57sffXeeNIIo1ESaNxIecAKZ+ViN2EzaII808IJrpkZZ4AciI3
Mfn6UXh/TWFv5vPfj1oY9r07DwXmq8nmRl/Swgk2tveoPhKfFHW3+ftdYRShz6P372ZqDtG3xPsg
3ZB5cxFCsHq1tprRGtJoYa6p9ls3tL6uXeKg0k2BLrc3MwAR+YJ7Hceoyg5kAA2vUI7cq8HfU4OI
5PyGwZ8dktFZVC9zYI9RaMrZPUrcelqKSxy6lfFpEzTHspnF/pFpjasjzOxHP4Bpvk9qEaHN667C
c7eGztVrvfHTL1tuFKoaziCxAB1OFcP0nPmTRgCYoFsj3ROp/aAbME6snaXjBKDesRwM0xHl38Dg
JolRANxm9GPXl84uZrYlgIgolxQx1sFNT+aeiAfkg6z/cDacxjiF28PlEoK37Xb9OxxUCXAF6ILa
OvuGqcpzb9Ffw6Trajr63bcafHGUVlpgH0eoUqs7nEkF1MaHnMPTn10axdzpytqewDiV/zlj+iUY
boBP/sxfP4KIJYEh9y9onZDqXnC/GOKwxXdnFHEkTX/lpbuNvhlopSP66xq64PN6JYIN0FN1nu5Y
ozCejMfPfy1dOHhAsAGS5QIQ9JoM2VneJwIyR/8SIKS0daDElQdB+J1/ywDn6woopKxAK7x+B7O6
Lk3uadhQjJ0zLs4lvIm2g/VkqV+g287RWZxqefc5dnzW1NlETfwTZG8oeXbnnjLFmH8qmBCyqiLP
450ZfhwdNeIbbeOC26s4zxz+pFRRdA3b6k4FZ3zip5G9UCC3gXeWdUnkzVLEiSqKa9MJUxCLnCkb
n0IBKLNqrTiMTs7xBalXmMrj9SwwXwVp006C89Gq8PeGuw9g8aA0ppeQvDeXIHUTrGVKBLRUIN7X
HrKgpqfwP6BbXeb/u/IEQ1uufXPGehQRaBfVueMCScXUjYWMlfq2X/L+A4rYgkWGKHoQkQDjWOEM
jR5zyqAsikxNp1osMe6eKU5OHS8kjbsUpKq2WqU5llRYmGK/lzfnp2tKh/jYzd3RXCO07S0t46Ax
KcRFKjT7GUDIlveu4N0PLAczlTl1oQCfzpMRjQ0s59IOArrSf+caLJDO8bhFIxCT9+ZK2DIjSh03
E+ofiRQg5FlfBGJOE9OgTIbJoDYvGvlscGb4d/jACugPXC2iUYMIz4ykwq5X2/noowEHXz8NrQVJ
OUinMukHiTtqZO/uGUqTHm1CwvFfb0SWQFFy+W80vgaIEcTLoxUFdWFj2Imf1G4YRZvrBiz0zWgX
ViYpUyrkn7bNupFF5buz0fwdnwhY3nrxxuTE4X41tzrEe1UxSILyw3vICr3SjPuK7lztzHBUxXKs
Bj5uwPK5kc4gUMOoflwSuNAIeLltuFTubEgat8EO8OaDD3yzXLqJE8bzO05hjg4XmYvOdPXwpYRk
ed3DZxIn9pX1PqbCa59vgTKq01RquLSYXmILyTML+a+IKvnd3Q3VFvrp5S7eQvnuzPxpQJmIStK6
eFQ9VrLCvvmx+cdvVIsenods3gtX9bGKb6x1bshTMsN55NsglImqS7ClbZ+X2TL9ly9ZzrYEIOta
brH/h47P8aXNYqXQYzx4e32UZVHJVm6qhTl1NTz2P3Byg/BiJWAt7mPLSvkt9tZpw2A6WyB59j+D
gO9Wk/6VaUTtvD0nqJWwR624/tr7aa5ytlAvZHUgqOS4lpeJSCedemai6ne3/ObiZGovHqmavsFb
V7TuI5Cxo8H9RwoJweD9NPQ9BdxuUz1AVOlrNVO6BYypsTGc++YK89ROaDkdHpDw2Bk+hPW+P/3p
0IZ61a6JAXKdtObTmh6ZQh9xKxdNDMMEKPy35r3JOWN/UHArYPE5h16VgPugHP8OyDB4x904DP6f
akXo9cIj/PZSv3/E4hTADimX+kofUkqy0URtaTUD7pNs0ZkF7NMjYC8HveIE/9inEUZTzZCP+d5u
z/W+9lfzFUks2O4yrDuBQDhpRTOvh42MxkxYVmlZWuF0jyjkxGcoV7E3xJly7BUkAkMvnYqbZSuf
Wt9U3k7zo10H4zud0PTEjV9PhfGsaDHcP6Om75qRZ5dJ1Iat+oWBnWWF0ke86jT8AhEz3RkpKgNq
Qt0rIuIItTaUhXIJYdC6myjTvKmrHwjM5f4nJW9EFvpAuvrrqLUYE5trtY0V3qExHUEfyOTPW+xo
R/sf3VBJZj+RmpVRJgT92Pujk/WpiVCRBj35Y+Ed+bHsb7/ew+t7f9a28RKoVnh5nZx+kxmMDbFu
Mg47YyC/OAPQNSyZkftuj8McZLHh/ey2UyrLt5tBKduv8A0tTRod9R+szdSNbU1USlx1rj9gXB6T
1gLxbGqZhhEqE/NsxNlc5qXgk232BB6rXbp42nTwWvJ+aZMMtdMuqnTtmBK48Lu4tAnI2Zyel1Vi
1Wn4MG2/Dd2E+OCkd8R+To5vy1VfrzcCecXAGqdPbbgow6+7PGnNIIjZ0hZmyqPpDlZepLxW2o7d
WdMv5lpi3r2kFjPs9dDpXoA1B5C5t/4CjYxRm8JeEiHZj8CyDAGUB0Scl00SMWeH7RTUJdFv6ZvF
0lYKXcCWeicWIshYXZbWFIsArH6gRBc3EE7BDdhhDdd8xbLWVtc/XXMnfvCX7IJIvGQKCfKxJLQX
EIwrDZZzAGQbgzyfl2argava1rA0Tw7DITbAneNzYsSdJ/2o5Ls+D+4Uukh5zyCeJS+r7ONWAycI
0mZxqZUnARB4jcA4s1Tn32Ve+kVDeuqPUewV2BG4PNJSdmMuowowZh3DNDBsG6uDF8nITEUJW4YE
KYpsWZfV5QtCK7ZdcjRtgE7cBmLH6AAv34lKEoxXLnpjFI+CdNdXe6OX5kUQB4IccXcMnlSWNi8o
TAYk92cJUEqJfu27ynyEXhkq5PpOjNtQboQbzkwCDqZLh2yArbqoN8KjahcFbrwr3OKsRHsFsE9i
1NdzFiDctcOysSJsdJ4pPRcLuRj1y2USeY1Z0W5MMHVSJp0Kt+47r72k6N22g2y/o8a8Pbn1PWTi
uIZ+7Du0U0m53z4OnjM9LwIEzXE+hJ0bVwPGBwmcHaCMfz7C9M0z0PyHhFdojsUmzqCr7NaiQT2Q
BbAOS83qIjjFss743zN+JdjT3HCp0su43J8UYbr4ChaJQ6+vGQ5/G4hAH1dk2Aa4VG3VOWiFUac/
6SWA3LOZVZ4ckVRt00BLUvEH1gbA1rKcNoef0UJp6RwBSorkgsCiYLlcTGZujZs+U31KIv+l8DWR
07u019x43GnBVLJd4Mu3H8ZYn9/W05BqBizq840RcppiUjDhQe++tEl+g2cOFonVTvrRudF36Xkm
Oc9HydGE9VvMVQp/5P4No0qQWWGeWIKG4BFPPY/Aihzzh8Nu+uIGQiigEBqfa8kBbhC0dHACeTmw
GHVFGOC7n4FWtojfHiRc+RfSLtI/mV7Q07BN3GWPPHphSmfhc1Q4CQv5cn/zVTQWqAjmorvN+rX3
qVPE80dYkD1l32y+uphBhLjruhdzz3hvYEwPXHCOADAVkJC7cWaiqNY6bkHWI5rkwKC4j6dgW2In
twzF6mIxn9cRIGR4V4AUH7lRbyVPc03yc2oopwuSSkU5KK67YRsIu4apMUDu+LlxoSdmQj/8TD/K
VJL+BUw1QUZgagu6TCU1Fz5v4HVmGCRvO7vb5eWAzG+aCY3tpgcjlkxBmjO6Lqkq7XjJdywfY0Xq
Ok9Th/sbDViKLs0PkTFBPMBSekPaR+PO0t38WqjdVvONDV+2sFfb+Gcy/tKzknqUFrcCWKvy9J64
1YMDH4VAqdFeZhPFEGLULTsayvE/uwgMhVE+Pxt6yWf/cY9TNfUXsEs7JvwzjJT15RhtOWikEJuJ
CckBdSJwotEJ8wBuuEmJ9UIwepBIG9bm5SAiRIurx+bz9DP9Ln438UuKfD9H341MyiEiSaqvnOZb
9k/8bGvmDNeS6W0AydOccY+gCRJGePhM/MVzah4mJh6uqzptkzCTgeV9PYWZH6BBhJ5kWLvIDund
mECKiFfub+cj6bDmC5f0iaWAAaIKehXdnZHpfjlJ/857TSh3/6CeYFuaJhhv1Np610vujFeiDSuk
fmTyImie2U6WWPwHBQPbwIq7l/tl1acYREonYO3X6tY8yarAVKB5PzipeM+4RbfHQFjjf7t6TDbb
xy4XYCeofMUInK8bnBRC7b81V62CkCqnVyGlE/VOiU8+SBymTgCAmG20eHcAyUjLIVUA65M0vPgY
4jNDBtjbCMOfGryYHx3W5Ghdw8DsVGCi4uat/wjzlsfaRvV41oDQV1GSNM/T7uGXfCLYZrxUvfym
mDLKroOsTpW1X3K0sBkBGgmoRKT7K5IvF9xUwMy3e7et808x23EchQRH8Lhc0TZVJ2LjlbI6ya6r
AtVRaYRKPxf8TnH5bxoMGofQ0supKpSDLkU1dI8GztA4uiFGr0UcmD03cFKwjtY3i/xyleackAf3
kGs+2atJ1M3FY56790XkSOV6nNar7SG0tAOd1WMjUuF5aPEGoD6+9ZbXnc0KmrjNI3A9U5NvTh6u
q/scPYxkKKL9qKzv/r8mR95yk+eMSuLCLQLwUNEVSW53VCzEkz85u//IG3Tb090At1Ux46ZX+w+P
IdTQ3eKbGASgSNTxyiNNvOhWBKSwSoXRZQ6aUslHysPceY8Ce3a9b96+K9WkECPXDEnyg2BeBH+t
88ZNv9+b6CVBs1utlJAlircasTZ0dEp0gx7uCtZRGD+atbK2Viy01C2o/mBWCyclEuUSpQsiMxLj
KeRNpS92w2lkpMvO4qjbuT97rlcv1XxSXuIjhgcslKRT02q4pLeL9fzFJopp29LIuj8Yb2nPo0MN
m1naEhFhBRKW91+yL+bH825tGFaiPGVSOVjInFPJh/t6oNVfmI7L5ymLxP2L2Ss9INwLZgir6Bge
phviDxA8YEwxL/d/s8lN5g7Ea8k3mk+vSb+nKR81bqsUsypSqwBSI/hpknyrWeX5o0CXavIlmKSW
bd41N2XaXZOJwPHG2kVzato5FjLQdwnZJJJW9gmmvcxlnx/JR04h/ksUzrhOwX4r0hqjPhFEkere
ZjxfdpDIDPEal52gBsrHhmx9T7HFhhN90hu2krSEqmcAbQvakz+0G/8zWzpFsDUs+Jq5tpKjUElA
mQ9LNkhomm2wql3S+g6IPXI7p/+h/oOU0Hw9FtcWpdWg4AgmMJFUnJB0e6qPM9N7lsXXTD76PiFS
yeLdkHawckDWc4FEJ1it/qPOddbm49LcC1YGbRQyHahS5dd70tgg9qH1yDgY3Qg3lpnHZoafnE4M
kxf7+UnRO0cLTbiotIf87RKO/a/rgJPvZKDiCKEEiBgB1VB1ZaBvfQhvau8MHcy6opaaq5RaGfOZ
Cg3hajIUqtikWMW1CMYekyI31Zd+3fE6sAB3+CUO9H3vDMxXr2WvhlGAd/oa5fdZxGZXa3W2CToV
DYFk6Z5UHskyC/gZk8j1bkYT16VLsz72AIRzR55ZQG0LEZYoFmD0+fxM5ymP1rgck1wdb9HVbDUz
b5g90pUwq4z6dFZkEvUXKA71FtVfz3ZYhlVY4OpzLcxCbKpeSlLk7YdzAvbnxXw9XNxzwoMZzg26
lfieHo9/Qf3stgK07ncYAwmogiNJZY8DF/Fgt90pK5//e7EcGjNQlAXP1hyhXVXJo8cB0u8/saKH
g27QOcfEoJLJvRayKIDoT2bmK/cvyYpi1RxxUlneVQdC5l3B4sUQbhjTDmWZ1OePPuAX+4MxmrHy
9rnbd+d6pNst65qZgUDtkeAdE4TdpOCdYBhATy1D3uQz5lZe1bMmOkocjxYOUhEHCU1yUb3o+cbb
45WkDoH78ES47QFDMyTvTCk4ZwCzWaF9g4R3ZzPEvWN3U67GBwFYBk8dvj9zixV28Dw8r/mY2Fhm
pdlXxBdquM0qsDBC9mXDQxZA0jselrnroAEjFCC2luG2yRbYM14nrc0sM/CQXLwi0Ff2TV0UfvI1
ghaRePSHlTKJPvqEE4Mnqrpe4hDPZ73u6++OquOreFoLTvZ9sJh25xc5ZoVW6CIv5a9gLf/3BfCu
6/nNH8JRet6Ann+u+ZpYDuCn+dig++nDEfDCGz/Jivd6ieXTZRnQzp6dFD3WmAOHIm/PgFz+b3su
WZ1zJIvvbcueEJzMrW+WKeHMHlkgx8fACm/R17H/Gl2mRauzKNAlKbHivEQ6ptBLy02OSijOjz7Q
7DOv1/HvXWAmqJ/TklGUVlZlA7d6tPTg1kVcVvZ9igZcomgmZuSHJ3ALvIKV8spfAeaVifkAA2ye
OfOBmkmd04e0xJaEtFXINlKAZlTaPvcgJsmI+FMw5UldwyPA8DnD4/lE375A6DjiUrJdXZQ15tkM
FMxOg2EYomSE7p6trcMfQmRXTJL3KcSoMJAOaaqmYB4WsJX/9UD6jAMm5mxnOLVKbei34pjYl0e/
JCLjSLyp36U9kNqRGjycVQH/NZDkID0Lf6xuO96AjgwPQG9HNfm5WwwyRpAdNki5F8OOfCO3oP5Y
5sF6E8BihmT4jVfvJG1Ynie2NqJUgUVeisllgOjw6jApgwECA8LFVhRFuO4Y0yOtoZF1Lnz/I3fD
250aHKTXIZUnRVXmxKqF1JuPZ3Za2+yV1nKX73BA3179zQtRTNNLRotDEGg9othgEUCKxS7xgpYE
hfyHzjvGsufjHr9o9u4ud/edwmDM5gwqafDI14gSa3DgDFG6pp3GJ+cIdOCnA07WQn0sK5pMtT2F
PEIjz+OJ+931+w39hyJ335/YTfRCR91NvYbXFQXCegYAJXd7dhLvIvqqj9/8wzQQY29Tix1OARzs
p3q6XswOJkAPbjaezCag8d/FBV1vZvFbWIMfpACalsntfKG0OWjIh6j/nXQ5NjW8h6vs8HglDG9G
a6uqvxOmNZ7EdjMJSTMeoJBIyFEWrudmkHc+ClEmpKjp4RKqqa6xON/HZxrswFmrY0eZk0CTvLkJ
HhkbMA5TF2s9MPuM4kgBtorc3kioJGbMBuOOVLYgyu9cPS56C6f7y1EXjqLDMKwkwsSq1SyB5n0P
RIziz9piFq+yntpIRUPWS1f7q1IjuWFfcJVwxtOgEFu9eXOlUDHSgUFXUnNCSHAsLJktJylaO03/
1VYF4q/0IYQrMS0VhgpFdxiweWS0Pn612mimRxSmBxG5XruWyUO8SwLJUAP/HEAzKAXj6uEOuzJy
9pncVuwsNunGHcpOMhMddzJNs68a0ncLVs4jozdZpweG32x6sxhauSJw8oJtyDk+gNnFQAjDF+1/
4Xp/PxxMON7ECAh3wwPYKDsGYcWpnWQKAni/czWxgYqwwXNjTBivU4PUwMDYxLDiItfZvKswZbtv
NkA+pslHHbd/SZqNxs718ILZPXZLdxxnsURZ2J86ZYJhsEnuMUKunB2gAPyX2AUBmqgzJysSDYhc
4qHA+M9/bDLoCW+sbUIqice2Reus0PZz7zOdIr1oIoALhNhnd9PsbFU3wzRbgXrlDMg9ftOk6sel
nLG2bv4HvLk2TRbcDfCcAhCdOtUQuBhfgqxyAkHitEv6WizDWPOBDMxoBIp4zVmhn+ZZEesIzJ9I
t9F+wZYrssKEXpB3R+HEsfJPCHcLt8GfhDNZKqC+f9l5Pi12ZvsEX8O1Xy9ESIeBdWi+NlYawT+F
/DEMC4zsMQJNAFSXALMNd5uf9iPE+KjqXy2FPOA5N7dBML+b16GTO1LpunQrnD0T0oDoh8Vy61hx
GmQQ9HPFHq2nQ+yMr6sLQ9TRNm7VwAIaPnSn367Fteh9hxtG7ztnYvyxZLAxUeZhFrnjeHn6uCZW
ijVVF54kOagVIeWlCCdygPcXIbB6Vt0lLT+7uqlbFprC0ps0SJLtRabvM83hMm3L7RYjCQc3asBb
3bbYnqDUUckSCJ1Gz31qxQmexB7kqaKYHovdYkjpFQ29YfOccCCv3AoKiUka2OmJURodGbs9XTUR
CXiVDiWeDdW6GK5yeqhdVs2E7Mw/b9FA+4y2c+gTofvST6Nc5Ck4msR/jnOciuO3ysFdJARku+SN
nMc+IUuvh7/Fjwyy4vQxb9dKBgbi2cZMZJq1+nUJQ3NXWttlM2u9BSAn9bqBBqCDlLw04ldtUC22
rklzCf68PqocqdCJEClk3m+gTxpzoHPdn2eI9g1fyIfLqqYZold5+cLOIEsmAf2DRSuRrBrsH5JI
p++L4dKCKkcCXQmmsyGExMM6tjRFLReDdNmVNjmHJBfnotKlg171ehFtt4ynG/dqsMYu8bhfIwrf
YtEthe/UNMoHJIjGM8NPdCYlfTpzIDcYeVHPmQiRvhl/pmJcW730fXTAMAB26mhGn7bhxyKcjvHk
+cNFzxxX4l3uJ/R82AxPCw4rY+DFHeIRurAJRAarB0X4ePLx5ZF5z+gLyqSUNKC2cEfgR1ktRtgy
Odb6FRlIJ052PeF7Dx2/Ug9xhh2J7699MS3poREHAW9eM9z/tFNQK9IzYBqpkAqTajiB85kOTK1s
DxHoVSTBsKJYZZxnMftrQXtlNwJGa3TxgjrHNlPTYofWXPttxcHwErzbk9ga9rWdNtpKc0sZqPND
e/Dc4AbKr63sFXb0B5aCFsmAxsPUOSsvpcXTxrjsCWcuNUVg1IqXH7sbmTu7VIlzzNvEzcW+8uqM
Xvezv3CieL82sQRtVcdiuy0GCNxDIKFMA9zt0FKlaLkyH9LUYa00x1DBDmY4+WomqnW+JFcexIei
sONjRqzwmucxx0qp4UkHmzYq3hJ2jQUSRylgMf0uC75SRd8GP04AZIv/izpmWA2rFLpAf6wV6Pz6
61bz7UwYjhAufZui3hbcsVBEIbcwvADmCTGL9ZaHX+Xy268v5KV2DgyojcuIeUteKsArl7x85594
OR2qYXHRsFeOHbdEnSs4bIdZixcck+XCCe7H8XSCouguskwqcr77L8w5trYXCf/H5h8a6KGLIVna
UUQokDCkoZbjtxmgMrNaOSAXClz27InafNgkjhE/BRwk91eiLotq+bV2iYwQuodbdCrn7OPieL1z
hKUQHawWZ6ImSohhePbnR67Jsa/4/EVjm0b84H7CDMlkOC4QMlkLx3pUzyCnbO1NNkYEe3RcD3fV
nMdJbsWg/OaqcprzS52V3w/7Gdzw7jxsseI/b/rKq+Tk/WkV0KzMLInR71ITyDN0FBB3tHv+y8GI
NGVcr74+5hOvVqX/RdwTO7mwrht+0xLb3JxnjNJ51++JxT/CAt223HpriTYAtRHx4ksh7h6+xDmx
eXqnlcrtC8NIWuLAlC9FLe6+VLY5A5S6zOY17hbwbQS+eAggig87R5E0C7fMzjDk5qvZ1OUBfy0x
XrtEGaa1JTiQCdlEaJXc1yApz3U5KMd5rBmYOROpHWpBMwLMFIUnuLGxxOaHKnTqiDWjGbB76QTH
UPO6ovYLSmx8Usl8l8abl1OzRPGx/epO+1rhfqI53jZrmkR3R5ZAadzBhQQq2sHdh8bFs9gAbTPS
bDzQsrZZhJX+N6Dz7K0e+AmU4XCmrF10p40QAvXf4rKhsQSyeixXCBKY6P+vYDy1NfPlbnCBL/Rn
gCGloBpVl8Cwn+7jArEuylu/ebHT4UztfSU5sGexUEbMffbFRNqFCzvWX4zTCHHjV1Larqzi6eFF
xHznTcqSmucN5jri9gamhwxSWW4Xhge0BTBOYXprg8h5mtcsy9CsZcenc6Gt5025iY57wDEnPycd
BDdmy+jrgzsFVgxD0ZcWwE3A8Gb5/FC9mzVPnC+gp58i2/RQvkeVSN4zu/41c0K3TWBM8mLGYXEl
H3PKsveBYWOy47SfDthQ24AxmeI6Lt8DCybMe3B+9nAFw5tc0J5GTzdf7A16hIVDztq511es4FL7
USK7kpAvjY9IGqnvAsrM+v7kGMHkKAsK6vDexNVHf6ta+jEq9/WCN3MoFT6Uj//AUKxqAihB7aT5
M/n8961TxQpRQlJsE1CCUEKWw7RfprQCZcYfZ0Cqyxs8l01hsldHTUDJ/5PRNU5zFx0/30le0+yY
0i7XKsvl+fjLc/OON1PKbEaF5BJxo9lStkFjhzYNr7kkpLrcnzCuROuq0U9F+qX4dmNg/0C/poOL
hxRiR/uv6tZAJ/9kqeOe2heF20vCWk2NOjAw/E447ARTxZoCWOLxEb3rV8JXDszsCVDMODZJ7/RU
yAwBBUCjURNNp/9iWgZcjyH12LRQMc1koH7JuA8xKbMbLz5FEnMNqBjzKZXgBAZg1yHeSObI3Lf7
0zVrNxbffsTUluqF8pp3cbOHnIXHyUu4dHz9MAn5KzHbAca8OjxdL9RGYlId99/OVBlnLsax+G8/
AIKXrtBxCEdnTqdgr3tQKnCPUFlb8vgweopvh//7zHOmGPW4XPMwfA0F866wZIBkzsDinlXm9hAJ
Yt1pD96y32V2J415zv8GJ+awK3osgVa2fM5+w2k3du54kevo9Yvd7A/i0Oq8jNgoSTuxfzzvTUwP
4+Wnf2deIsx5XChCYHckofQIUqKP0mdFFTnvkwzG4HD2Rz/Ewgi2HVSbCJrzJB0MHGcQxC93k/eC
cUhgEFHN9nt/QWC/7TAwnIHc1HrVi5zXU8WamFbEd4zxCH6CAtE9i2R/gj6rgbGM3uctSGwTfmKi
ZYv80TO+xuodJhQPDlVmJ2El7Voq5/6/IaPP9q/P2bJiWZEeLFYk8bFRvNqku4q5p77FZlo2yNLK
mpNr7AJNF0/n1nU/N9aEuqU67pbgZ5xFZ3JwtRCp3Khv9WvXT3/T76wCOzui+RJ8dOOGvKCMYrsB
tueFq5prULqc9QGaNrjavBgRFz4ESUFbRw4Kaoh3rW/pjeGnHPwIwRysaJZNOuA2njDhjt8KNYHn
Muf2zwrhTWe0mxZ0RS39lbl9f8b5KTZMmM0lWJWMe9kJIEsjvnku76riFGNrW5jSlF0ZN+Gb9/j1
U0YolzRRjqixEjxFju0Vjtn3fpdpgm1jLtS1lG8kxLQuOmkYfKlcd6Vs5/ECBKivwx+3CQfroeyB
SUMGhvSi4Ab/7e2DCoOr0s+aM7CCwJZ6Q0DMwJraayAA6tZcU+cx6WgkYXIQJXDnALszDepFHqaI
LKnenWSDubllXxS7p0Vv5uXwBX4La/WYlGbsDq7JlPJ2d7OVeg+gVuN6Ht32SvjdSDDevmkxKP1c
hdqsUsCuT7NeEUbKlkYcmD4W53YmGgpcWZEToHZ6Zh/XeotkShqAuL3JT7ryrKykbywE34Q1lC+F
MzjP/YbqYRfG9L+jeT1oTZzV/pk/NDqmdypAGzLgr61iEkcKf/V7EM0VoXEt8SWF/vLoyT6NRJfC
JsHLaoXhKESE6TTDnRGDNiU/6EmIaz+8dpTu6nhmAP48icmjpXAVRYbToupiXHSGsZjXdi2guFeX
AwcwvOmD7g3Uctpe5PSSiZXs24na6QtB0UosUWq8/fnI4A3f5otVI4elzfpO+Qmc0iGvBJ9Pko+r
31x1zOt01vKDgp+NP3pyZed3Sbra0y3KBMSH2oCpML+ufO9Y4sRqGwaMIPEH3p3VxV0uI9Gne6Ax
9kwXZOottAYFZUDHe6Ocd0mRjwR52F+SYOnuQyOoJZIGKTqKJ3Rs7CAqtdl4HdoqhWXYm9EIobAx
iRXayG+RGQMCcHiW5hefAXDunKcCpBQ/gY1xT6JO3cn4RHH8cFltDW6oUP6xx4ejdYpYm1ux5i9Q
mS1vWjfi+LlCMNmvY8suB867A8UuTnqhUYfxzZlPHiBI58teOsQtenhvgsk+MDFr9qIHp3yiLVY0
v+jZ+VKTwp6vej9sjBwx4hcfWPjeNVBNtF93yxCq96HEOdr1VuOWMPxVXkxsItnNbo4bneLgnnPH
sxh7jbra2f9Sn+p5xDJbuhNsh3iupBHLm7CLidYkEP2J/GSPJXUi/zdoQpTcP9LPvCFiDGzWvdoZ
awnL6bQxO+8tp8Iu4BhSK4sUO068p3+7tTEKn0meWytC9O0albFiKKr+UjbihYu27O3Db3pO2hPb
NtzNyRK4dBdOM107VIgSlWiOgZ4Rsz2STqL3phELByKWnZOPEfmeaP3Ty92WCZYzt8aerr61ESGb
itKeavvcJpOm9Sj4dtuAEYh3dA5gAwQ1gB8BltY9Dj18gwV6EgsbgczOP8l5eoah3h+apYDstCeX
cKQGPJKhpV/fiqnz9LtQP3e6YDOnGUosJQI51dGJyaGmKWgeARjjNh04bRFPi6xcz7lMWHeaI9c+
5KzhYuwRdKI4fQ4yfdMgwCCoZFVYazeI1c855Ekb0Ex0bwXW/M5Jp0R6dNfb2puPpWCkGZtiHTDZ
SI8gqB3pXEnBT5avqY55XbYV8kmTPQeUTAQmhqmHO+Uh4GWguLZHNAoFEfJtYKbQTbnao+YLwczj
NwG4AEfvRuOhXd18WelR+9aoQT0l+fTuVo0Tfqr1I9bgMy8Ezo1c7Tix/j3tpahTbBUzYwUoFrHM
TNn3jhzrAVk0UT3SYtqfE+VJ+gG073ObfAD2ORMR2kBjdNMQvKOjH+fMXF3NNHKiEqMFOvKJZyKu
Uu/+KXZZSEo2p5hyzyRz3zZKts4eKGgsI6L2cS4z1uQmaasuQW1c7GvybjidVw2xLM5lxp8ung4u
NNAzwd9kbew2FXExpd3s383+q1RRxZkMO3MHj2RARUlsQMcoY5tERKiPtRWY2PXxz1bd+RZLrUCz
ED/kKgJMUtIZ8zDYcPs1wPoHYb9n/Ez883CzBdrOnBax+mWuexe2J9dob/cTFU+dKn100zEKV67S
TDEQv10XWjqqIpGGTaCXzKxPKXGTe+H0vlegt35t6fnfUHw5yIc8oZ0duC9rVI60/U55f2Eqj8dx
qH2sZAyNHCBTIR/x8YTJOXvsJ877TkJbue/0J13xgiGBO3NnoNXOW8aOGdIamIp8YLknVXK26WKq
vWSkNF65FIcKPDNxllNuUjKdnmb4jvjW8PsNB2I6zah2wheq49AWhEWjJ6FgUDXs/a9Pr+ekcU+k
PlG5S78iI8vtKdWF5+FL+fIIyikDv+Ra5+FbtEtbi4LskPf8s+cloVAsQrt4C/QMtgCT08YCtWdM
0jUWPI0vGOrYgg9D5dtNADz4WXf2DwSWeTFuNIpnBYhbTQLkESdOHZx3CoWyXvpaDoNDqBt7zhLx
6ThdfExa4ndxwO0Xgm1SYff+4buhYw2VkGCyuW9aCwmKd+DBx2NKKYwcJ6aJXE505nMYUPB1MCiH
MqylEUcoJaRJv+Ltjfrv4iieEBmiOr42jXg8E7RyYL7vj/Ue0NJEhu+gh9ORgmIROC80kyvNa9hl
LLS4ZwG+ZwKGYfixKcczHOM2Za7pP1E80UVl7NJ+bdcX5vmnTLhG4Hf9G7ekRemdnuIO8WpC0y7u
cQvt/i7riFToNKn14VVeL/Z33iJ+JeHaH+G0FHsQckv++T3gfrg3Mh1w09JXhMCcog9JmIKRO/VI
0wa2BjRpjyFC9F4yGgHxRi5SXJ1T0Quw2XqhPpFlDFcU2Wpau18a1pAC1qXGXraL4XTK7XBMbQy3
2vjc3khNnT38RjvGQ6fbEn94eLb+pj3ZY/kzplrU7VciiBboVlmkcRMjBY1C6VwUcknC2XF0RktT
2V+9tfXBfKH1CFgPUU9UIZhFaEhE4bi1u2wtrOj7lAhtmb3H6n+qSaJ2iKtFNVuss8Sa0/swkked
tX8yyI4OHIzLojUTcz1ttOaKcP0sCQbZNZzVk3YZ2w4WlbBpv+wCjRz32Z9TOz4608T3GB/nbqV6
AHr96/bG0WB6yTUFZGfFbCFmQnAbMBFGICU7stEX4zmeqUQJOFof32e3LKugakJQBfi0fWcrRnzz
lnwxwvdm7TIZIKwAUdLUU7yhdWiGqn4AguE8geb/D8z29DICjws5ycd6Q7CpVCEQln/WwVqsXOLv
/1YfXPnZYErKikX8es0mAdiG2NVxF1xcPjbkaiz8ivuCUSNGsU8hWtcKZYyN/hMWx64YJ87K+CEm
WHHzRPByOq8S0XJk1eCfwg/96NtzGXy0ZVwCSwK0CTz1kbVe7/WdZN3JzIbXqYsgTtES0mazuRho
Q0aYVaA15o4oF3egT+gYUkJ1Ws+17Uau22NlASX2Y4zzmn5x7plCZsmF954hEjjpE687iNTTyS1e
N83m5yMfBGTsA9BrLL/bYk7fxNVOTZoxeb4GBuzlbvNl4mGtNtceF2kjFmrmywl4oqJr/5s/ciOM
Ypd6WR18V62Ox3eCrU0OV9TE4WmQCbSYSR3uKdhbUWhXc8ceZlxZ6LpJ+i41kfa0Bbt3rBKK9jlB
d1VuQAIrEdxAaHUzmblORnYgDr/pusjJ4s8WyAjyFYdeQejKO+o7/g0LK0keSEQ89TabBwHd5KPF
xvU2qMUC7RoT2vH3+578rjn0kKFNpO1hyORzl8AJL/iJ2lnPoF1ACrnr+Ib5IStlKc8LPlKowEtC
Q82UHZZAY3XgWY6UNOqcXKij2QFyMsQdQnFp0GMYm4POInv/hywAsGSe4HBKVGeAazca92WKTVB6
nc+OVTFtkdaFpwzBkWAyYwQVi7SsW+xIKup6CIczboDBuN1pK9Quxu/pHFg2f6Imih91kzDNDlgh
lOwmVy4hnAp2W7pgFtJstV2pclhNNnW6XFNXlMUpjpL0KwjBGWOgV7/wR7E1UOU2H/CC8hBKXmPi
sPBR/cvD2WQxh8+ocNbfP0/ihN/vWMq33aXmRxOJPsLrBjuw0+I6LzixUd9mhw9no6kLnBxumSUX
UJu3twXI/7CDBfecgDRB/aZgwTThc3x/DLjcdvC+fUfusc7h++WQTNxiv0eW89owoqXAR9XwPhzU
9Lv77ts2BF5KwhTNLSLMfl+duq6fcZUGBdI3783e2xXlYOjeGnIvARR2QOhpbJDFATXBF7oi/g2D
+SINZE3ZM83pgIFFV4t9iHMIL66u+pZ+5J3DOJDJfZQ4Oe+0tjtVYMSemGnZscHahAz2+6W3icGf
rKN52pPMPNKQ5lf4urjADZR6ONtDjMx1NEXxWZ3l7vwnEiBeGR/QvisAReQW65M92I+0kXfObhjN
hFecLsYRayw7fpF/d7DUkgIn1mUB5BNxVg8M6BmGPWpJ0Z3yYZHQKINnjTCyKcFgsPswKJs2ZYn9
TUpj2nRZqWqEqTVW/46tfBhRpj03r5N6GeAepNxLoZ5RseSVhs2t6kZ7BDh4g32AmOba/r+P8nIR
BchPhT8iyY31HEi8/xhnCm2sIxngWyLxBG4xJnYAbByH0tnLY1VzY9KrrqjpY6UMRHQim+bfS+oj
4BbLheClCPGDlCG5ryHQqBvSMpculCdVhfZYTrzPHRmheivEQ/PmTkKNN7ahkEEyDIyZXs0RxfB9
NbURuTe1pW2xez2Cdf+2SbTDrRpSc/CTvsu+m6vW1sjlol2jpEIFn9qlatqCMT8TopJak/BMn29Q
Aw7Hr045+RLtOvl5RUfeQLlNdzNag+2CB7Z9SJt7qKIgLndnkg/8szNHn8PkcxmXnsSSqzttUoKX
wkGAOECBPFP8TcjOKzU0wdCDy2cScc51KgA/R0SUlMGhevuZ88lstwE9wU1edBGxbdzmi9X/ZgOP
l5u9/3fu6LMqd1PlZjjenquXw5gkKRWvKPY4F5b6HQqskK4Cb3KjfuD4C78vje2RtWS9QN8lKiKy
YJOArOu1R7IBbWxstvixAcglRfBJ9nBNzg54yPOen4znHQakycCUr8ig040OcraOX8ZJ/j/S3Eml
ITUpa5uoI2pOqwDMY9N91rVxNu/PmW6VIz3D8RkPImQnalgLNjPAupg706lRE+2E8b3H0lvWcveG
xEVbSzuK2xFCM/HacJEJEdOl27AtbXhFjacXa3ra738as3Q7AW46SwVOX1q0i3N4WUgBZnOaCgh/
lWm0UnKFyKz5Qe21cakezmps+0BAxy3E7bOX4c+6o4j5tJPHZr0xA2pLrfJkfbRgawiga7KZNW9m
qsJrI58kGeVYnVtbB0/sdoACAlSDF19Zfq1vd7vWV/CSFXAAwyLOQ26ZLyAzOXuXaAwCc/tTOzqy
8I1ke8IB3v1F5tDNYsYBmwtxY3fZKFbwwGDeDQZjkvLUQY9Ag6eyPoPn8yzpNUn3ltA4i1X4UKQk
tlQPhQNyXI+QZXFrRG6kEIZnu1+oADtLIB+EWZiqj15/3NgCyiYuYkWeLnXHqrtyjZhcD2iimr36
kCVUk6Z8AiApS6/4KFEFsIQL2XH01ZNTO+wPTfKm99yYFyoYUUgpoB7HLUI011oN6efq3rPlv8DK
2MFuMDLIT+CzLLNCcqvimCJ9gUzalPZbvOAauUbfDcAj8IuVY4hMnYMtzKwbvSgj2QPDTn18tZS3
nDjBREyn6D/7k6kJE4XIQZvigKb6Vzk0Cjhy5dlw7S3i4HfBnfoQJu3FiqTLpLjoz7FWebpanUie
ktBGXI51IkYlOH4GCWYXy169bYRruS4+X63ptdAyhBlmwWKLx8bqS3sQid71UuqI3AwxE4V4cjNo
y/GN9Ce4Vk84QRt/HIdniAqeFuYWUPkKdYRa5O0XTtByv8mChr66kU4Lz5QXydZiM1VoFJxiOuMP
e+yXM+hzGp5GDoV6wPJ01d0Zc63r8BRuwWjDicv4nCYuxOYRL9XgzNnROQFpHZJdUs7TRb8PvlVR
6/b/CeNgyRzibLdqCvFpTeEktLvNni5Mifi/WjTWe3Enac4BYAbyd/7Q1xN/7gIrvCyf+fuNVnE2
gDs4CzLrma6qzLADYeEELvU6CHImo3VMLZALoYd2QpszwTKzpBYF/q8TLi4+xIm1G8CdMPjex5QA
Qk/uSprr2UmgKHCox5ittlYiMLBnlt+ct/9gIzRzug16azQHZlk0DwR3nRltOZECKOuoDV3n2Xc/
FQfbNoU7qc86H4fGAb/163RM0POxQFf6ttXk6HWMN6dPtqDQbr1kRerXvsDY6DUI+oq461SMWwPo
PdLqaCsXyZQmiIdqj+Y1e7iZc+xg3hjPnzKBZ6AIiYx5qfzSSjbmMuBhp1RbAKW6WnejjjvL2wXj
BWV6XvpiiUMM/JYJGIc5AiTVr/cvywM0UQ/pqF+CAR19cubdRHp0q2ihll7vNnx3hsqcAoVC+PMg
f5ROBf4jUlE0NNA7R2dBID9NpKIUHXGmnjKtiZbqdYF4UpIDxG6L4JKi9AdFkgwShe3BDAottvPx
MRGa9hNvOmKPGNejaj3AxL7VVC2lDZCV1lozRiU/acAWIJ9xl9ua9Z4zYCxDweEpOwGRf1DVLGrj
R4xej1KKGhXlLVeah7CMk28tXq/gC5wwRXoxg7N+SO9Jdd8G4wve5yG+nsG7xEKLkCkDtXTf5fiz
gJ5Rd4U5yPUytcUeZanaxviuWTRd+vuVQa6ksa18rLqLwL27psxc2+NbPhZgzlj+3JZuu2hWpaD8
7OQpI+plArC/wka1vUeWktFGXx6bDxFOSfpdxXTFXCcau/VfakldOupE8xOOGUsFjcMZwtOJAxIy
3ftaMX9jIaeI5keTGjGzL3+H4h9tapxj4BeJ79TqC9BBTDDWX9n1J9KgkWEn42d6ZlHft2PMUWxF
MKWCw2aW89zOGslOlQ3uT0GBLt10/aVciusnDrM9n+1ouO51ofdCjmJr7zDzXTgRrY4sRNPkcJMF
h7fPrBQqpFJ/OHuN+PO8C4Vbkd8gAWqzkGbF4vxF/gQl5I1txBvk0UXFZhuHwxJ/kYL4WC+vaNjf
yUquh27U9ZPhpyqOX8D0DOeBXsWMFF3UJgQyvNVbDpthaFEj20Zaa1pkEoCX5blEMOtxuGM9eFpm
n5bCxf5g2QVW3vYJaO0rZOJ888hiWZQbrIvtvJNUj6cgCC7Nc3GvPYCi2OObx7i0++42T/giSui9
s0dqlm7LW06Qa3A7N5OyhhtS0Y6nVUlgQ/qez30NwK7WdSdNGDKxqUq6i2GjUWxU+qGrewVYNa/0
pFj3Lbxkr1K+I1GnE9YmQeQl6oq8n8z7kOa89FweXEv6fs16QmkkL0Ut3GRLO2iG4toTFYNIVPGR
GIvj/AsCKIWA+Lchoh6RI52kiShZ1lJQDyTF73ImOb3+tOJ4aLxlXcPV5Z9X6pU8ME0Z+K2cVvig
/X/92Y8NtwKgCH9XvknJ2BlN3kRz/wkIB70ZN+ZsNSqb3YV9Q08DXpIB1s0dtHvVRmPObAATMrKc
EvnAqZtLvdlSQeHpaVWPxuXJ/IPj0D10h47V8e8FkdmDgoyiRV7lbs8BA/Y/BQrsfHXMcGCrvP3W
zStZxelYtlEta6FskT7iUjzu3kNmTXS3cvCUie2nUJUxVAHQjH6DwACuveD/hFJay0Blk2sYnxdu
5kp0MzlXOW3BFEWrka45m+na0IYmeMa9TPHUDfQDHNQVoMUM+LocMmEt4ILxcS1uTfqGL/bxItXR
nqaeoTQWREz9s+r6YDIPDuSAuCQfnbLfeBpeRsVyUBXFBY7JpfEgA4DjLIGrZk++VLbp5EjadMUv
VXguPdYwwvnZeTDZG5aQLmLV9KooR9VuNjdO+phy8J21cdKtkRMW5HbNZszBrEY7KUTO2o03Jiiu
kP8ZWojmjq37OhC28gGSMZI2l6UcPj76aevhX1+aMFMtIyLmajDFQ/Mf6j/GZDPnZbhd4XFozj01
OQrLPbk8ZD55HOyjvr3u3fzbC6aL2Cz4fZd0zf02gKpk8q0oJi5igKvuOwdONw3jLwRpFL3XoaGo
bfpk2PcNOaE5gxQ/ZffyTKHs4W5/ANKvjrh6rMRZ0sDVuIR6X33KoBLuC3TGEzqw6N4yGIhR3M/x
wDFAUEG6wHL601lGmd/z295uGj2tFGUQ2ckH570P9iaz5B3LH8WBHZeqbnrIe68syo/LByyYGdzi
C52iMR6y99z8rE7buL6P2Na1ow+O2eT/HDw0QYvTdRR5BsKLVgrMXTuf0RvM6ps0wk7+NuGvzOPK
NPEP8kPGZNJeyb7UqTs0/2dq9nvmxlSzDeizWgRG9QhDfGTe7nGnj9CVvyma/4wjRn4IQXNRZujz
xs1ur1YkgIswD+h9qPuxDzKId1NP80ZvlnKsLUX/u/pyqR3VKM4zbsOEDgc+Od02HlFDYxyUMZDh
wxmSdS5dRzuANhhi3gjYe5nCE3TWhyrJZYJJtFf37SZPEeQQH0bcxMuT0vUlGHdyol07G5rnXXhN
/qQdje5Gx7URvE2RrDAIaUczGInJbH9SqiXVw2XTVCFDT/a2cRNM1cXrrKGDksPyVjmyTdLYl9rM
h5z73aXRox54oUK5LHqB2OUkgSl5VdlyTyGKfpXti2TQdLDuuw00tYwRcnPlMjl9ofrfGf7nmqEJ
yf/IKJwp5Ddq/FVi3FjIHBKAF4YPceXa6+0B9YnRCtPXZV1Yb1o/nk7JWciOq34Ra1a+kAWb56iz
pIX5FhU3sI3Irw8Dq87gGmqXQCGX9OYJIxBJ8ZlHssOCgTeBV0VR4FVV0uNINSAFJJeP+OQYDD6u
HDLdLqx+lYBRQDeK+Byt56QpzmtWrD7aQ104sw/7Ntldi5+oJSzkMr3BhEElkWVmuQPGoIMYN21B
xbPVDoWRr2mU44zzO+fVfLb73tgV3zYrQWkxe9Yxm39wvt+aDUZuLsiIiJ4Ma2oWl/+9NLRPjEvt
5FAR5JJpej2WJmXm2vemNSOmMNyky/fAbGQ+NVTRyMze6L/5xq2CeD2VTKbfWkCx6/oBWEhbdkoY
c54quDAkqWwqRcedDex5ZrUbXcPVHlo/eEia4GZzGgbdkv3+KGLsKQ1byPB1BM38lm9Mr/XMrRMK
ZuRkFjm2tAVofhTK1PUS8vhVvnERXelg37P2xPXM7PI0SxnRcr41woN7x0FxmsKt7NsYCoUb7FVU
ZqAJIGGfz7QC2DRA4rtARQKC3mB7KjfWTUAPdibEy1NHgcytIeQKhDMbhMR44KPVedjZ9I/rdi3/
fEtAY6WHjB5o3W6cEkZICUMHq7IOaoQ2pM0LA5pcS1lNkgd0iC/flJrPZV4BYtPlKCrhjbS4Ym3L
DznLNyOp/M5231tBH5Ok3hTVx3kIxvSen/YbkKD7FfjJh6QAxipuxso3JemdKXs4ebxAmMGSZf8p
VrN2UakMSmB93MCY4B/CTwSBWB2UcNtMe46ePX78jmjWQsEDIucaZqS9URNvozitWDRW6xzg4MRL
rvMqfP+GmGeO8HdBXVg5kbDHnNGEcYXgIayFBpsAtmHSZugQxG4VULgxvIbkPVXr308sXkh2XlPv
byjo+P4VXRGoKT1RABg/9/FD7q0XSuJxTNkjNWqcXYsjRd1G35sFp/BrUoiWetuBt9OAgJz18IxU
CYFHWhpDjDRjOozWHCj8VwUViN/dPEMz0ZDyQCrCcBuknm8QQc7M167gQuvAGwLgribxYycJSbHT
PsAppmZoXUAZq29ajTi8dtOEEAfJhv6chc/Ql3+cKHBeTHPKo6WaLHqfcWFeJUX5DSasDEqeVyuK
URqtbnEtb9CZmm3EwpU3HR6e1wpLD9GncqjnpBq1+NtQxG+d3sp1LkdR43mWM8J/jLocVkYDQpwO
+lI6rcxZIxWu+Et6Yuf1nBu8qjNyByAP61ZoX9EDQim9XNMRJSYLvPV1CliTFX+8C2nMeufOWWKn
7+beP8fZvGumg/YUpc2N5NTT7igyobFrufapxTU+GWfmV9lr/ul7AvAvleJJitXKFs9vKYvZQ46w
1o2DwCdVx8N/tuzKa49bdWNZ5EGNf0OcAgn3JxT1mAFxEO1hEZPwzcdsUY8HtzDDURnqdqhUGreQ
/bELXGnw+R17MAMwLHpTnbvq7Q0AVJht0be019l69mm+FO7q/JGzGVryDpvJWaL7LZVA6xEgf5u9
nDMG0kb+lQ8VeRDLwufGo+21SXxpeytPj6fr8h/1ihiEnS3NYdlRC3ThxAe093XITMLV7Vfuhf/c
OC5kdfho0G46zw9MnA5TP6Cd3f/oZAXZGkxZOCO/cw2/tcuRjWKcmnhaEb6LHagnP17FQ0R072QY
4gT+hTbjYG7avHy4fpyqp1ZDayXEwWMErPotVGPuwFgun1rZIgRDPmqGehaKuHWoHFnVn1DzLNTH
cXwT+HzITjtWu74ulmdSYpLpAXYpS+zjErIeKISF5RPMGU+R6W2wFSmQdVaIpAnBFhHRzQzSTa5l
iUnNHsU1NCCN0uAbuVBWkH5mfqg9dIEtLhFsUOUvblSyZEFEKgJawrElezjyJPGpe4oSJ6AHMgqz
i7iKmESS5d8XQe2+duE+Kucx3CNPHxzX6nXU5OpLPYnkgUsPBM8T8At9d5IeGu0kjh/a5u3fkVJK
h/kdycCJAgGpSuMgJxzxcjH/KjkZuv4nbSf8rkvzg14yfek4ImsAaxOXoDAKON7YqSLRiAVfuYsb
MiJvbdR3a0A0e1hL4EJLydlozjC0Nk9jrLLa448ErIhEc7KRjgZpKMrey+J7/H27RrmHsB07e8/T
0Y9s60Hz8iR62TS297Urs2fN2h7/6oVcHdVI+hshtP4OMVvqe6ZRMeLbzfI2syIdyC/YUkE1Ue23
ozbd3tbwOhBvurolqeCK4kGjr4BjZG9wA9qIoYwXi3czWj9PZtRLRkgsmTNBeatXRX9KqElnA/v6
Nm8Fd2+3+qLzTG5vbqYc9d48kqwMNWOKYmPHDgyYulWAUI02B6EOdXnLUm6yleg7/gVa50Elq5Qg
gotSvlaTb/wjgPPXrtVVoVNh8k103ZPcS9kNedvqaLmQQPXRR+VgVD0aCc9pn5NJXtfN+JX7ek2g
57K77XdefUpCG2Qo1dqn+dXTke9KCeeGWvxEf0HXR2rLe+5kOq7/WAGWjufIL6K0RalpojLQsO5g
qU7R9vUqSrtCGgl2yndhCtOjRjUYATIouMURNRbj1pIWd6YeNxvuRsYJRZwFcoDnI8yyBj625bu7
FkdBwKR2KUW9ymYfJPT2kVoGfsjHa+tJPnJnbX/yf+/QBGIkVazIVWrzt85X3RBDaWOv+5TUFgWu
ubnI9WJ6TEsVyIMZoXPCQT8yhGyc4uAj43uGBNUAEBPZ1VMTgWCcXCA1q2Zb8LBo/UHObQaBRY8W
uQAKhfhzXcQG8bkBFheP2rH2wwBYO9z+96qH7zqc6L6j8des9ltpO57su8A4VF5toomQs4JZQs6W
4S7cdfSnkOKkerus8uZRQ9yw4NdvHgiOZOr2PIS2Y5zJcvAdAvmCLhHp4QHbSw9kxVZ8g7xkiKuC
47bagviA7uJRhheRBNR65szX4NFpjHR5iWxtc07QEIDF+0j+xH5sv5Zdfdm0wupdRwz1X/EJ5YdT
9tq/Ze816SU61Tm+KHOmc6LeJrUA03m8T1KA7eNiUmzqNszJeQ+9C8rS5NNg3X8yqw1RX+oS5rcL
1eKccw5SX2ifxCp1NGtF4Nc8R/ENXN3euRyriWVm91y+nchrVuzUJcB0NVJUDh9pBgqm2y+BzhbA
svgQT0eapa/mer/hpJULw6gTAWU9X1gE6XRH4hOnuLhSLs11agVg9ZvF0xuTKMv4uFJopEWVkX9h
yWqhFbLpNRiBiws90dbG/H6hbFHP8IIWKzj+Vt+1qVzW3EtQxbkg/1Tvy5PTuCiI9Z+D6u86+goU
2P+o9SaWWytsluW8ldv8Dbk9lpk+QGJ0fc/27wpnMPCBfhFXlR3sDW8ED4MlphamKLHx+5Yri2HL
hB2uY3qG0MVXtpXWM0g2L1zg53N4f3pG2F3ipK2XapVxJ7BcDKEcqAwVDawyRlGyryBpC8ZU3hcE
gcCcG0+jMCoXQywN8/F91zK9QUgwNesBNhatN5f1DP6Rg++9bAPiwQ1kDaKmMC6/RdeCVGlPDJqZ
iI6WOxczWiWQH+h1RYfAQUQiH4FaakpLXlCk6+AOQ7dvxbWXN3zCitCADjvyCkyglWm/CKDgl+F1
o5r2BrqLXygh1IP919tbRTpzvNIG9PcQhCudUEAbPI6zVsoH5qrJ430Jg5/4xeBqL+hLjDeKyuIK
esaPk5D/3G3YmREFREP2zF6jPzq4K4K70lWJ1jqPNJb/zr7BP2t7NVqGNq9qdSpODz11Mu5wkTMm
bqwkvtPko7WlnFH4vMaGHXakUnEamlsrx2H7em8dwvBxWPad7wwzJOlWYqEOzozg2JkVtZdmTMEp
Vt9A+tRdhOnvmlJRxRc5G+4WytfOqxuSvMquPaDoPyf10N0F1VmSFZ9TwBPmiMuxE4Cbv829LgH8
LxNv3enDwygrNC3pCQuDYkIMgXQpN0vtRf8APUelvY8Ik5XQNtKzwMMXQ/OIMnelBd5VTeDhbXuU
/GOF0qZcmVHFWK5s0lQMPyFKC00MRar5Ovkxm69wqLc35WF30Q6Zbo0YDj17jJZHJEP/9MlS7Sbn
G3WH/M8u6eHfHq0m/65YSja3gYziP6l6YBCKi5i+9z3UocFMgxWZ2i+8Dmp3OdbrJdpjD421LY1Y
Gc62NRkZK44qI2qzvkiuSCZ3boij0ZfWLiQwlZ8P4oPvNjkKqE9xbtMasyMneFPfd7qxJMb5aBAz
qpTSU4B1sbX2IQYIfwm/UnVz69Bu/WiW5nX6JahG41okGMtOi2CUO2KiOgixLqcAP3zUoLMSf7d3
PMWhwhj/6tmyunjDai6MPWNaZtCp4TUhalFwWw+k/6EzHXgk0OrwiVriHAoLZmB+cm9kVfowbGnB
h9r7w6uhaDjoo0ulOHDo21L/rH5So1yKyS/AFNwIElCN+is+ghY71g0eP0A2R+QSTFB5rMf6qUdZ
ajRM+YPUqTiaeqtbnYaWAO6z1+tg13ZuAtyChluMMRyJ/GiYX53qqYPx7UatF3llURzIFvi+sQ8h
1AfO2nl3klG6F9KxAd6PBDpUlaTon0z1JOZptOUOuudlleAVMp0abcAeXtAsoIANKX1qv8EoHEJI
5sfbGQmxyfjMyh5nuypzTP1YZPHP/PpCDk2O8nkGfZKvI7z9n6WfmTNZ2oatMOvvghlT97DWgmxn
4aL4YxGxK7+YN08FhyQLnZ7fmDK3vfMk5prgWF3GGaaBuTpTRuE9yCZJjB2QhSD5THDI5ZxItqs6
dyABRD1ECHYTYgxqvkvJVH/0nyB/HW4ffadAwTjaJo6oR0nLVeGE5HMtRN58o0lvZlK8PANjaJ8X
rbcinvWY1eEyf8TfFZ73quvLkTmD/SoI/pvbp8WZPPBkbU7O1g/DRH3w+QTaLnXsrJUt3AJIuShX
iKGO1vi538+v3Kyye9IbWCcZpRuaK/RUhePe8ttbkbkHm+OBLO9DjHoGuywcc5PVpNk9J9aHQniS
DHEIps9V8J61x8caws1gcpoipTGw7A7HC/e2VpO76ExjNNcwiGVwGp0GayGolJmF+XTd45w0KwHm
cYMzWzGNP744JSuFSNCUMRnDR8uJBBVEMXRMmZMvxQWy3Uq4pn0RtOCilISHmR9LncZcb33vPxTK
trrjXJSRRaUbHe7+0FSsBTB0TpQKQJdFJTcI1vLjppGh7VaUqWfPJsvhMLniX7/pcYx2rNyDqpur
JHWdhWmAzkgwJoEKiJi1sxSHM2G7VPvwIp+Se1jzqQ5L3/63x9N5KXJaYPL+oImTOYHHe2Qmiw6F
l/MPfWRyHc/JhC1apdIV/dZOuDHb7AZ55wZtdzE8O2Ayn9JRjmTUmC5tusvYCv0OyegE8kWjbxdv
RJ8tM0EG9FYjk3XuHdNfps/Amzn9EZWxgn06Fluol1QESMwfrNqdw50/4diyPt5LSwnKzKPnr66s
K1CzNnr712MSYtcXtdl4ZYxueAYloIP2XWWcuF6g/zdsXCWLYbdnbyqp2g+lJiaRO5RDU+jq997U
TVgRUsUwSID1oFlQDhZphllPQEJFZ/xCkxWPkEnBD/WyY1kHO1HfFmBY/c3IB6gTQFgsTSGUY/v1
cGLJ/2SLyk+z1WwAC9AS63Xnko1xpSxiSEmgS2gWqDx0LHIvb8qeqn9KXopdrfZC8OOGSrF7qp1T
KOjvyEsde7M345wEdE5gJLc1oMPUgCJAR98SbpvfzGU2hx8UpxdQ60/u/BNNaPJ+oejpXAwB9k7X
Z4QG8d9RTtKjpj0myQ4J5ejECIxErtGY7kux8TbcfL48h/TIGsAXHorvHElt7+mEgDzjD190mfq0
8JkRr8gr7l2yNsRWE2uhDm+mzTk8eHy2bV3cBEZCSLk7hUBrKnYS5vKszR1GVbRxLCGZK84SxEsV
xK/W4lrB/OgHkP/vUs9b0aOtN2ys33z5kvhSD+cFTJzFDbborrQ7eE0K6AttJB/hIgp3Ha+4NyVr
ePJuveW5OlCmApGXZBpr4xgIIFvb+odf++c+Y7ewJqtlW18n3WUlveJnTiiAHuGN99AaXJ3dvCTl
rNp3Ycd3LwK24nlHcpDtoyCcT0wPh6NW6hREmEwUi1SlfM82ku00KPaOHJKnTvChHCFY6MhUemlc
9Yl5xnwZ5R9ESG6J4zfpFsv7hypsXHliD+9/k57XalR2LHIaDLBuly1zCIG/ILFi0rN/ahpJFBGb
/nuUDd2/yQrjPeidf1Fg5k3TOjQUukYetWFOpVzKkGDKIQil9xJNHANcffJG5EWVF1MAZPSsk4ZR
eFKm8V01A2Z9u/xTTyiMuy+kXiqC4NrhpCtyPspC8WBGKSPaDDyOxnGik0B+Dd5fmzO060ntxvx6
G09yfm278wHCJbrfarBPpOfbVqCLJw4j/OdHZ88daF7ZrxPxDi7qOlTuXAiIVcSS+QXwdKtr6vaS
HooOYoj2KsDYGSGLdGWR4X5T8aQ+TzS9z3HSJT5btqE51cttOok2qMslRhLXJRo544DJ4OpMl/TQ
Yk6CyJ+eiVM2Yusck3Y05sBao6i0OofFc5C+mCTpz4AdGxbCx+mmn9RErjoG1cZ8S8HQqhegVbP8
C0mwPYK4IU7MLE9qsocG4JBP01kYZ3nGRHgzCCLckBvxLf2nr+hSX4cciId3BUFv4O8KCJYFVuhj
lELoDg2QG+IetfD7alE1iNvc09CPCmYw+p038Jnob6dMpm2TjmGNv+PqPOlKy4fZIoKYiyBCDoyw
FMNZ1qLfcQaAL6QrEzRDnf2ua8kitr1L3mk0fMgueHxODSVgVpMUcHr3OKMhTQYpOIEbhZ2Zi4bP
Q3V7u6ll3XnAL8wh/amyvZNsAD8kIpGpLsWSbFNplLZj4eK06CXHpI1tlSxVTh4hZyQBf6kHQpsv
F+3S39o7zymZE+g3E/J6p6+0WkYTAwlJYT0sEL/UeogcU5mTXQq784916/wHzwN+Y+xntLQ5E0z7
7lSa403OQKrzU4ey8ZKobO2YCDu3cbFl6ToFgZDsRyMJGq7LpAHb7WU3hrbn5qowxuKzG9SFWGcp
keTho8mWDxCjU9rMs2x7Xk1iN8gyUmFVEO7cO0o31kJfw/CvVp9xagv0XbEMyDr9Ho5Qb95RF0u2
iVSCd1vDrKDJ0GkjN/Pu3Z6WYeHuGE1um824r6dXThdU24x5XdAuOBhOQfO1RtcL7SzQgKWwfMOW
nuGVj8FC5iNHv1lPy1WEuXHhBv/+bcYhhJRpDSNKcMojTT5Q6g6R+lG/cl0iBfcnCWAnQ1RPJ5mS
TLbooW++YVI5XS933HAbi/H3zIrKdilZQa8qfB/OXoEw+6srAQOHUD5+GrRfg+zSO0It1SbwbvTL
c+gAySpfhPtw0eLSPtIO2iW+0FUhgdtX91fHXza3P0ZZJmFByVGVEjmljlx9SkFYShEQP8zeIkXu
X7c/Q3cYJklEYYDw2jL1VtkRXmSNj/2yxvr6qkDSGEoVnB2LZGhzm/TkRfb6hZhrGWd3rwY3tMLd
GdG0QbHp308Z5+F4EYjzF7W7UkQWRGC3PvwUnnPpf+LTBthXNAJyhtcfP/SZVHYCxFEt98CViqlg
Jvkc2kPT/v0aSv5KoMZ6nMcwj2X3ZWOJzz+4G7p0l6x5ousF0tuReNYq+/ywf9Pg8DAtpgw0ra2l
vSBqCffreazIJ7lkpM5ZnWLaFrWiwE5cx5L+jTh81p7Q1sp4XHSC9uo4a1kEzVaK3vDn4s32tifC
QBmB9YSAy8wiC/Nhg6Jvcz93FTQ5zSLoZDPGuC6Xaj5eiVtHTNV2Uw38Dy+TDflv1++uhR3Fstzt
CCVMXlRR3d5tK1QgybL3JhsEKJ0Ao8NdBhrYZ9cPs1dULJM/sSEgTFVdFnOpi2t9iUc+QnEKmMXl
GHOGXUD625kCUtLCK6Jx38Oqcg191IpFu/Q3v2tNx7bwE1oOjPp8P7zBkS9SOljqiCTkxADk3EAR
Cqa9rWEmWyBeID5dzTZPLhSktLL2lBc3yQCJfSJCldby/2HfvbrEqmcKKo9P+LiLXlbYpGVXJ81T
boKFxi3SDqpbICgi+5ObG47H03GCodNf3ve2TjMz7f8yfIbRztATmktXSSn4z4bZcLOv0YRkZkDF
8I8u8rTiMta+U4EbHfnz1aNzq6pDI1OsS3dM/vI5Mq8C1HE4EtsAwNBvZOZBoSEa2sgzPVxnZX2+
WOy2YQ7R07JLE+8ZCOCBPGgX7LSHeG67SOY7hiecrJOgQdOciHcx34+uxgPIbEnY49Y2rm8LgJ7J
vYaRlTnh0oea910w4KRNe4N2K4GLDdyTKSxOlbmw8FjdYA/qElBsqhd/zTaYXKGYPyJ3Mq5TrlPo
tXox1pxwl/AhPptzYlcVzezsbPYo4OkUytxHZ1vm+2irpi/8r7F4ZoSwqzacVWRPpnHYCETa1guY
RAG0f6NOUOSh3XHaZHi6tg6xBqoMsnZgOUFNiQrk4GK9PKIBBx46WWskIzLvmcyZCKvG6dqPvTvW
dgvPya/6q8KwzcBz67emVSgung+vi/9r3pIrzsQ0Y/nzwm9Js7+5Sm0NKF+FC0OIZ03XefebSDjL
tfx0SiGlF4FWb5Md5zws3kJJ3c3X4DQsvZnNUZApEkOKhnXB++6QMPOCGSA2OO+Y/S74oB3jse6n
dg7ER75/0LwkEJjfs2ujyDSNkxoOHP/uOd7LglNH6xaFtVZCMBGDLO3ZYG7dbwXhvbHH3EJ3/6nq
PjemGTZJHCUOp47Audke+LNUO+YpJiCEaHcdmq16sd/hwHi2n1bJZ7Oeuy938oZuma/mz7UtfXKL
bNFKe3LdWG8tY0Ai09cEzVX5EhziL3QDcoCkC6CWd0ROHIGCwa8EAxwe7kbp+VtR3s8aejIu4w5t
iyxOx4vG7F+vvd6uND8p7cpcu4/md/8C0RsvhL48gxyVE9CPdOPSp1WbJJFEJREei31A1GxB2MTQ
0WsSWmprCspQxW/1bfeoTj1qYsU51MCWRCJn4Or6TF5nqoP3EUj0JfFpREw4BRLAoW03BuizdH1h
smZVgVrnImnVMt54y7Mgcd66m2BdjmJVPqPggpMX3ratAxKs5EzalX3KAa+yso0ExkCfUTudKnPO
W+WgW3E1aVs4uGRBnO63zepeKiDhKbg7xQvkInievY1B2nKDArxmfg8uXNBv4UAcoZsirSgONPp1
AY+3AvkUa+dkhuoWYWOtCa7in0xe44o4qxOCja0e+G5wPRSffLIC9ZXdDzclaTnArMWOWTBdVx0w
lk1lCrhnh6qzEdHTX3O5V+qQgdM6JrT9zLRlDcPmd4Dw8zNCwvi5GczGwJDi+VyVxomN0vSLqmSK
OLJhBJxWL3XrwPwzVx5NCrnKleWhuaIJanMyQBNLKAIJYFgVTADy0yRG89FC93JGNW3Hsirh8+pq
GhN6FfAu+vx3tzamjWa2d5Ez4xj2LofYeopTOg3tEtCP+mhCrewi6RYRQO0xR8vzrY34wNUcSU/k
uG4rFSx2nbRITqPfk7rWejsA0Rw9YSsmWxvAfURTLxW6qxRnl7+tt0ZIWJe4KfdiADnqEXpdpHk7
8C5R1yjtO+DHQte5jT5eGX2EYVUjRtyE8H2UCQVSWJ+nL6VFyl81myWEhwEZ/Y48JX6bNLREN+Io
1PWi8izaWiRv9dhs7jpQzlDFJh8B4GYIAK5cqp5zeCdCVrQsiYzr7WPNAsioQDwZat6ioOWK1UCD
CX/RGKDf7u0b9/nNmHPg/XqgNJSBXOY58N9lr9+5XdHlj/TL6CLVPqEweZwsPxZELHcWgqB3Rc+N
cpLn2puM+ZLIsOcA0e5WPfzhhIr7R66DqlDxbhXDvnIhvdV4VvP2oiHqwdezKBaAGVwbegYUXlxB
H/JOaVBsC4w+evG4XlKzqhl8qkh6LX9XV/tNisXG11ddNehYEPvlCUGbZCkwAbohnRENnI6/A1aL
YcgZ+7eRXmmz2Q76evSNZ/ps/nlQoCdlIRwqmTH3p56lOddXIV8iB3J0sq2nYTHO6/u74Wr6mkCO
GCI/jQV+O68CwgKabNEJTPdOVjoBs9L6UozWfZQ+VoYuL0WQ7yaRHe7kKLgppqSZT2Jw06L62zA5
idQ8YINbPAhbQXWMBF6P0pMRNZpW3Lvh42Ahz4omDVVgzbhrafNPA6lWm4Fm/iOGAONJjKuwuE1l
+qd7VCKXKHBWAFxBDjO2N1eMnEBvGPgCDCULBOn8GB8nTUrpQw8C0Hw5fOJ71LAGrzHzmYc6YUtk
cjc0fFRwFtM+AETIQVtZQph5KVyJhi+q+WzOaTmy0fc43Z47mtb9jvyonoYNFfsdxIg7qg1NtlS7
vmOPDY5f467/4c0odluLAsQZ+ENwUtPwsTYb+yh3G5gUbyV411ILr4uV0VitBELK6DwrHPxCLW6Z
EH1ahM6hKW3E03+aUlmuY1iymbH+Z+WB7rqMgC4FOyciOM/e2ObOuxylAWB3RNb64EZHJkoe2TCa
dOVQOfVoZIz+RPD+kwg+k7WRMxmWGIT9e0eEwkhIAAhizXojQ4hTme2Cqoaq9dybENbLFTxpSdk4
/5YKIgTxQxxXKH390hgYDw09KF2WaTfS0VU0Tox8tZGaAgwNgF8XJR45VgXtwyxWxq/q9dI/dCI5
58QMbUuv1otfp8qiTgB1NQz4ATlJcuh+2qsPQWEMuiPCpzuc8XYLWdGi7mdpV29rYodeogbV6g3p
6gWvYgW7swh+g5wRKCCsi4aYB4m5tWtwIH84BgTsFZwX5iOVDTK/pFASMI/l61PZ0iTzEDsNaabN
ounnc063hcgbm887MicKyn7lvDzJhe1C9gPvs1D84+hwmuCnhmqBBQVxqBkAAzxHtHgmWHf0FSm8
tYtCvJczKIM4ydOpQDTGgaW+QyvDNqzeWTTllNvrXAyVOmZ9ss6viSNla06KbdzUrxJk4b1DFNgn
sMsQ15ei0utF42ZEUkVX4Bg5pXPitSfuVI18qQ5iZVnfXArR1UW3MAO4q4BxjImsjc67Ut5qdXfl
MRGBvRv2L8RZ08NzUVm2tnBsSGvBFMFMktUIv6XRb+n7R4Hc9v/mjvmi86eDCMOT82MF06MR/zV/
j6wtbgBCnLMkrcG48DxSY9P71SWrjvNyq8bXmGQlBF637Qxt3c+d1qj/hTE7dM+4D9WJzo9nX0C6
QZvPn3DhVLKJVHSNtia+sW6qVmA7R4OVJlO7E/N7drDORn2qtbwp1kl3hI5FMDspBYDPJWQ1rAaI
n9XuY5/IZGP/c+7TAzZDrsXm/qyMJ2aTsknJFM2P0KDSR42FAv9N1ivxka4l46P0e0qD8aGCGfBp
H1DPIOffLQj6HKAMT9j3iQqDjWr9h0nKjim7/7iaCl+Ol9VPyJQ/8xSQ+UsayiOhW+Jbw4BAIpwv
uiMIh5h79smsH2/unN9fO6uUCmbUHdJ+AmbSn0LbyyfSNC/2k2CcNPG2mHiaU5sNGStL988yjZjJ
+/7pMZXTSD/LQ4kcHWiUQpLDaHWEs8N5t3S3Awak3nbvvqkUcuManf2i9R2t4zXRQRkmmJ4k5Lt6
NDzRJrAc/MqEa/fQ2E7Cue+FgtLnv2IBx92SrxXKqXrZtZwqNpSLMt/sXvYFViTJtRFuK2kfCHLa
UPvpsyCpME9EwzGzucF4R1Zj8gxYedgklVwa6Zr3bqQC5AiSIkr4dq/QbATaUyc2UP8i71NooyeO
HNriswxt+tzKNXVST/G9+v5IUsnaW/HQLLV7nIR+Ap65VnA9GRdgGknmW/8NUj4izhxEJBqG/j37
6HuYWuq04+N+qmnoOsrO9/ni0ywD+P8qtzIYbfMSaLdMFWWBZqw4LMZDYmc2BTI/uPaeuMYrz0T+
zzhwzdN3Ghdzu1u7Zh3Tu8ITe2cdP1EbO13BQ9TMi3E/H3FgA2QKT6ubHSM3HB1IcJsjfwGgZvGX
mQ0qke8JZnMeF0dn76gxGeDGQPZAzfd+VOdrLWgYqd0sslWZgBYRhlnm/5qHpZQWn0ZL9vPYqJo1
54JlLPZAxuENktC6HUj76uzuI2o0UFFgZJV5uNJWaCnrhR6S4FUZfSi4JRYg8oBBOdv0d2dyQssl
70lEbUuAazhvisSuzuWRILPpWhBkUQzJOsH3boGpRzS4I/g04pPpWw7eR1N5ZyDtzHO0DgFMjI+2
o9gXVEaC04JU3wU8IL0v/yMkeLOJ7lvkct0PidpJvKQi6REdxZcBqVZ55eln7K6oT8EGFDHJhTPq
eiPFjMkeuPB2oB+aHY2ixpYY9/Sk18qhN5fG5erW6xRUTdWfWuX81aLImmy6Et9FQ9cW3eQxYvka
Rpl72Sd18lfIIs2hbPqie1OB/pGTDcFviCAUnvJkSxiIYc8/8eOUz4CS1M6gfm5cUMduPhwvidlJ
uoNOcw5l7GbCrc4gNKeihmGjvvC6fBcYi4vpgB8dARgaB86czk/n8WabtkTDSx2qSyjfZmIN7HBb
hV+dNyfzO6utqAx7gBxALPOCoPvEIhvsUWkgIqVMdFUGZT7bOXttHLPJvYe+63/5dTfM+ZfnG8ak
UGw/+aRpAfV5yiBxSGSwbDRQn58u+gR8FQU4BIcSWBORrKgE5h4xfc4Ypx82qBsEonXVwsa8L+Ji
REaY/+fFwOvswu/MXoVnVff18i+dHe9RoCit/rk73+cL2tBqw601Z5sVyFqtXFPy/CP8Sjgeap0g
yuR3mo2GLwCu1M9GBQ9gCo4PE/hl8Cfv5dCtUzocW2kNPumK7wqDGm7vxhUofCa2hm4ebiQq2XzM
uQN6deVUomTjyDl3Ws7HC/d9Za72OEq0i3mdfcn872pQWXyGpcp1Z/iBoAN2tRzZf06M66PDBbuV
IBktNsg4nRt4jCRA4MoXNfR7gyO1OuehU2pW5hE1tL9TVattMoccWuR4TO3xuzYhqgeL7jtENyoy
+xyPabRnrMPAgk8/fOwTVw2nrb0cH0J1hoWDGuhReyz290sb+yU39j4jDX5z+6Iy9pLv0PrmsR2X
hvVuxX0yjQg/qfDE4VfXKthSkdhYhyHTLL77tsX3IFs8UrjU26gprs1485TAcri/gak7rPdXZbFA
ssWdEGCe1q9lhf5jQbKHeBLpmA4wHhmnIJNky8oddmhr/W/3NooQCEB29fa5xbHpkrSTL5lrzXnV
ffBYEcFhgkz39ltxsQLgkXcDM1USfo/xtZxeWJiV6UM42Ns5H+FcnQn7CBSVxHVbv9VJ7YVcleGw
maZnJG33DKtUJ+MZNixE2qMfgDU0r/drE4hIQW57pphkb2oaympwAaeD0LAd8w+x7lHQ86jbKJqp
SOUYhQgDHSwDuMnV75S7GMJTPuGcnyA5sXyNr3LAi/uanEmC+U3Fwfu6RhQPK15QZBvaUN5dQQGY
ejonED6YBf/Im6NXnIheUAmHGhI7yJD43xa/U6jwL6RRyhAOPj3ZV1HHT8JozrGYkXGMjiiCSxbr
ZJv674PUh3nzBjXqUS9W68zPU497LueshOTAd4Vab3QrePcM2gdL9UfYaU5PlOpMHP4Jji4ySL/P
I/EY8yEMOpzDNSgyZKQKqUlvxvZLXWUVmBKaGYbsuuASGfdr2zFesGZmFzFaY7kPmcVZncKTbq8J
oinpqv3LQX9SptJJClWlmMkP0d1TRbCFOy37fewxKkPAUBuV+b8Lq95uC01CjuGZ66wr1JXL0Q1X
YNuzSTNx6Ldrw67wgvJapr750E5KRbu4tQs1O4hzS6VPoWXIT9MhqgsbVl3OJu2uf7HWQdQoacj/
oK0JhW10PsIXz7nHSpeHpXHSGNtKiGXoAiRWVcld0tz8eoZ5SC07DfMih9sp9GI+j7KcLydpNghG
N4xu3XIVGy1f9QzUgMtPLCG5MvAE2xQTfktjpBKVtaYtURnZZKUHUpPnPuh4MXjdp6/f5aF73+sF
rTUhKVW6AUUbzvk6r6nmSOkYlsDKSbcWJNKmGIQ+PGg4tLzXulKWJ8QMXXpIcx4uksdpLOqwd5d3
nApOUnlMwReCglz3L6Us0LvANZJnpisXE+KEbZyXCBYu6ZiSJ+nj3brtyEm35DDRuul20p0ND+W1
QhX79a5JFCGW4iOBtcEwG0fCxD3ZTSifPAxNJ7EYghTiNKS391eJvkwMCR9z42bTobqQ/aYlitT8
t8lWy5ubGcl/1/FWKiWKNYAJzbaxAdDaJiezfkh0uxZuqa9gWg8csIuGdAu8BL83NxRC88cZYVzj
qTgU/qpxMzhWpcR47IBPas/KNag67Z6AODIFCD3XZ1JZ/3OSWpkFdsCbX09nKBFrPqXnPIKRQ687
7O2zM/lBEcnIFT2vxk52Yvcl2MWXiWIzvrRxo/v0eHCGZ0QzWexb6R7unR5mvrJLrARf6tPwUh+e
YV5ZdZju7rPQFLClEygYJb7KJCxzNxpqQXjbpa5sETaP88Gt702VcWmo/l55oZfO5jQ4/QckuP4R
/34decQfmBTHI9iEdZf8fFNZYo7NY7EIdCeT0i6XuvYq1bOUHnzZXXFiYjAFLS9VCkmQTetF/wQd
bmhj8PBBqGGVPquGxPZJJqwn8jaY6vNDuWY0aLAF9nq0JBl2/z6iy7oxd6CJs+w80ywWlSt4VMqU
/Hz8TrbG8Q1jek9SnOSjtBsRhhVbcdDylAMyO3R91+5OXdaG8l/KzmWd1dmvw1z3aUenlv+BZZ6g
zowF3OrprTz1z95oUpSnCqTsOg0wDwPQ1DqUjPe4z2VlhNcEzs58nsg+TccyPbahEsC8immRyKdM
h1Dk+UMV1bfiBXD+wmKcbihQU3ypaZUQdgKeOEWyRE7w/NELkLWzaW9huEhU7KMDYbzAani4xuPo
2zhg/zhnpU5hVVbeVzvMsB6V8O4jbX2FD0/JIhG+wlcDTWRctQ8JH/fTKzuQzVn+BcDgqd8Gdem2
mBos0tuZ+0+NV3G3OEapkvJVDh3g1iAoUTvPP92vj69Agn2N0QNvgJt93S4tY79dJgERfzOKmT1/
FtFEaORfXDScr+CZ/wI1Bcjc9oofvW/mERjn8jMdtM41towpp62WM78ItKwhPrHm3nmc0zar0hYw
pyLN+s7FuX/bRNFKz07+5+EpeTsOlXQyrLrD2TdnQgRA7Pb3ATGjk16x2oU9KlWTu4NiH8Fg1CLj
T1AxPn1DfSq4qjIVUPAYdQubZJNQo44bmXKyqu+0Z/CuV1OsMekjXU6oKD+x2eQ6t2Gg7h0xW3/u
lYKJtXoYXj+9Vu4PHtkxYVj4xLvmNf8aFDmmE7kzZvaBxnfhikYCk0t5MD2D93Jv9tbbxty5+Yau
0D7//Si6JEzDec5Z6sf46XXusD3jmSIuYxQAK2401ObM1Sw64AAiWtcOvYVJjpELtpW6iWp4o2Qg
5ojly6JrxUlMD1LDeAKO9VlhR+nM4bSh7Um79aTkDRaClFdYNYB00yHPbTAArhTzpWXzOA+zmMKi
t0CVMVAR4Whn2/S0hEBxu0p5iPD8C5EYfAZOjTcQ64V3+g6JyIl5MDQvF1nW0zTyUt/iqapnBa+v
SG2J9NXzHqM2WnekyE3v57MjDVAqMfAG+7ghjClTLGvG2Z/PKc6pBfHrp4l60UNTBQATk58D/xot
NrCUep+lJfJOaZiFSZbvCwN3biHvYT6BWDP2jK4cvIvYyXXTeS+Mwr1+DSNZkLilVlm0BGdxODHr
V+0uM8k09ZdGGmPXElIyFKnaIrBeGzGQ1Od7z0qNImk0tBMaUMGRjGjpSPIS0hc4Yg1z8PYaVEij
VZpyKb6BZOV7qbJb7zvUDbBsAqzuKl6cJIy9EC+4tObZ6mMtGRBrBgzuql4M4I7hTEoGddR47lkP
MPrpV4k9P+zajdpUFemr5qm2vLkGwKF6tsfowYJcsYgsuMbzgblXYWY8WUSVy851SOL9D/7ObQua
2+V3CxRPLVchZzo8Fs9Jt3y7rebIGQyQgoxY+heBHEpv5R5oP6eVaIMhO4vXZMRPgvYk3vKGHFnT
ofbxT51gskPZP1pz9DhpB5+sw5VExYCQS1sm44N7aPbcA0zhP7SHXS5Dhof0dMBoTsh1KGLrRogD
mqMUDNpExAc9QkYV0enEc7uc/wb+wRdA4Qf3qL9KjMxWvwGzotxunVS+5kU1aj7KQA1GmGgnAFZX
YI32qoWHAuIcoisdNR19naGbtE9jpeBRLy/4146N/SS4k4StNOINdIgc7tDq49CvKL3Nvp04WNR5
kFMunMeE5a0wnY8a9tX1JJLDn7RUPVmfOs2RMbZdekBiHKywxTXBqCM5Y5PpDNgjpehZjvlYjc7i
eGh9smH/Vulb6Y2bq6HwvqGGn/XsOa9teythSci9ezVZSRcQDRFPaR+JaOUyZvfDdOLTx1joHPDI
G6ezn4n9dvdmoMhR49YmHjhN0BMd3lWqbW4cgCWU34BbFmIaeDSHqSGuE6zRpcf9OGSG8pb6vxA7
P4SBoyILdVqcAb9utB+sbLNi/20pgkLjsc+d3pCdxuuJvYI9AaK+pb9MDeOiADikEEiG2XclFbtD
czIJDE7LwW70O0gKCYIY0341T/6SC/11DA+tvg4Dtwr/O49NIlPrZAmUXdkufEHPkEZEq2Bnrpbo
dclYnqkq5LKmJYTdK0vVuWXJztkhXM3ouJ6ZNdEXgKkBtMoZbOkqIGeKyGHuX8QzmcmLi1FjKbrv
BWWpSt7kL8ccPKiu4FaeZR5bruhNWOzf3cSgtSRjog/VYRwO6i1v7VJJgcP83wa11JHRcrZJ5r/m
kNLpI2UNPqbkWSsYxeAMfukYPSN84suKH4QRjeHw97kON7J5nzDraXBpjvQyJJK6lJ3TBLe03GxH
b2CwTVzrVVk915OTfSKdNDlf+wtWkJV2dLDnk+75OQpteGKFs59kNbMaLsVpRS0p35HjhWYQKIoC
CLhSZy7ymXj5lWwX8tfaZubWWdLlFurSFTJf9iJLin3qBSetc81pLu8DNXE3mCJOp1uxIfHStYLd
GJKDt3EXjT7ILZ0ojbxP7/dIc2Mk+a68KO6ZqKPF7+SVunZhz+DSf4rLLhz11bnCLwPfMHIYyV22
rwCpVLOl+Vh0Pjn7N9AF13idTB2ZR9jA5DKTaag0XNpOY1XHz8BqgfKKqwUBe/xEE5xRnizzsMPI
VdTw1TbLrAC8YtiA4wxQstNZvzJK2VdL/Ud5oV/s/FOZYxhbZ94/GCeK4OpBw0GLEdL96pP0FY4M
+8jncRKK/9MFRNB9OnOrH0MPlW7b8AmRzusXf5wEcqMdBRlvWRjOXdUTp77aNFYZBN5TJ/HuQN/l
eakgC9KrLm46iypZJq2I21f4r8amTJPV695ovdle2CDuFjvESO+fwei6TKJOvbYHsRoGtN6eCpdp
yK7AveFIm4fxhbN+LGUxP3VLNMTtiXnZFsqOwCVVEL7CE6BZJQ20vicPoVXgTneQRjVPv0yVy9N2
TZ/Rdo82WffHQBF3/hJFkzpFK+rBdveEpUTCQOZ4tmTGGBOHLEeSRpod3sqt+gAu5+rUZ76WvP/p
QHcAF7ZU0hgf20VmviQuMO0VGANxMraa3AMojGeGeTHsUg66HumbU00b+Mgm2zRGL217NSi2+yxx
U68AYtdXnzM2P/ujATEt5IqP+agkPQiGfStn56fsGOVpQx/3J45XpiAb8F12KrWzWqJWK1pZv9/E
65bMFM6A9GH5Z3vHtRORVk6V1Xk+/uvUM1Mbt3nAkS43BIBjcAljoMAGoMBVBfZYmzh0nzE4jJ1a
m3UIsqZRbPjZXCqfBr5DQha+Q0Ha2edABxZi8Cq4KJHDzfrTx675p0R7yOYd888l7xuAUm9CzCL5
gTKzISZ3VcxT+ydbUAenRZ2YZ6FyiTGukFXHfCyjfDgpBcgfrtA4jGdUcB0ZIAKObg9zYbZpzSzu
dPzyc9/6UCL6xSZAofhmgVunfTgm3e694hzEFYK69S+KaojM3S4KkoWM+CXZEfVOIoxQ6P5o1O58
UH8V0eIN/jnMzY17pYKm3FYdTR05JSzkRa0nUkejMQnlAv1JoUsOfMm4I2wqa2ZFLPVz5+/UHxsf
6jZvuqPN4lBOXPx8phjhL+RiIuwYhnstXWEY7nyONcsUqqrw75M0/KKbXEbPW5Y8kxAvichhLemH
7KIbOrkCbf/CsmvrEJvdHlWje7VATIhmcEZFixOW17gFmb8Qz0b06qmthNnaklPLAbbWOyvam2sS
sSXykefHwH80Eeq0j8pMdzWE9ZoNqNTy+E/EwRr6PBGs2R2jzsJAqP+hWePJrxJGptlJ+eyB9tQ4
yTvIW3MD8LZEFh/kqoYd8tYNHDqkX5rjETPkXkvQBIB+fWYFv/ZbsukiIqBUgOzD+5PIwsOYty/7
CSOb7OjW/YWNDCB3rovzSdoKuDxG/3rcfKDJPDIDDkJoU6iPXS99YrGFCnEV8UBc8x3eAfG4ln5f
dGDi2isqfLujzUdSrB6c0XUeMLmqLbyR86FbAZbQFMExRnWQj3CHwpIQLFZFxS5zB3mHib6pfxL6
6or/dCcCNXz87nUUr/Na40IiTrnLFjNfrw8G8BA3cvDqUgVaxQxLueQ9wJrvibW1wclnhASfzdBD
9/JX7mtNewnMK6hknOlbKE70s50N7liqXalh1zVNc5eIM+/dFclKNWG5/UtC4hQrMCSOvrOnvx+w
xkhRhQjuFb550mlwSRNwARpN8HrDyaJDmVBYbeV60xCJCqRqaTN8iQRh4JLGM6ngdZkEToD9BVhH
ohVpaqjWUuokh6qbZy3TZqaA0qkA8KEKJmvQFCNsvaGk7GqlNmdxVaRLSGz6SekMJAWjS8o2Qzxy
Q3BQAF3NUGPIotKOPYPdPhxpyYHs3RC54U2biboELfo7Clj7uvXCr7u+PAMwSMIlthxUSisPcaK7
7f0A2B0WtX5udu2d1cp4Nd+8LurOyNkjuyc9mBJHJg7fgZ7mc6RTiGj+oKi3/HaJ64syPP9Fp4BX
qyL0fW/axNIuGRxeNifZj78zXFuUxgIbflNe9lWEifoyfE4vKUAdTNuIa2btJq/RxjZugNdR4M/l
3CbR72Ib5+9+C44Xg2OJAgDCMe/+Bm2rfOB24exapDoaM2SzK3oNDY3H9wTQjG85vg3bID9qYklQ
rpe7YDxEGqm5MtCkxb1C4Zkap8SO1NpFUQmGRDqoAQoDA1lMoN3xdHjc6/OpP1fdgphpzThSeOUZ
Km3MAzJG3mRoV5U5oXbkiXO6ZLstVldVwBSjIuBRdX4M0iAT8AH4+2UkS2panOKii8kFL9kpxg5x
hTyG6zbL5mtnx0SwQKubiu6GtMDx3D+UXL0CEVLs8qnXi93NrZMfQCDLBOUK0YWesXmsj9Mad8V2
SHvXQJCGoQ2AlSMnVKTpTxOAv8/iH+xAMiEM07LaF43MFmmd7GOzK834l3tgzSFSj+p7KzNLTYE2
d+4wN90aPm73aYlb7aR39glYbjbZDfn7NKc5Ire/jcn3noxaz4EdI2WZ0Auc7ufDFsOQWlw2ZkJk
014G9MtbaI74UZ5ot5C+Yv8xs5+OzC84q8kELnGErsu4EI8ySoU4PFM9CBcGaVvtWd/Q6pOPP6BA
lWgXaFOdOPwhnBABR/oQ8YWGoV8EYCO199ZXb4/K0gZtdn+oGM/um4HtrEyPhoCDWT8oRtYQnU3J
bX0tBSv3VzeksUB3RGHwPQ/0ajnaKxaWNTS8NlnRNH+M0aB/v8LFQ7DkTkwvfM/tBoCPGsi5AGa5
Oq5Vz21/M5dIQ8FRKIdby8ONX03h7xGGBRprig/RzwL8YySjjjAwj7MWDnAX+it02KVuwvI80Fay
QYu+kz6QbhDK6JYXScgluAuxBbE2GFBdIkCGaIrVKY5PSb0MtNTZRs2dKg03J7WR7thyiLNDnoQD
PBGQhSNkN1RHOYdtsvsXCwn12PrB3mxWeJXZAcUuWhdH8xzT8KABoJ79GAAmBEUsZc9KI39aUTXh
t+s4OmH+suh0rU0sKFgwqAtoWhoBXbZqTRFO/Gq3fMsw1RBb7bm7UB6+Eo3RlsiGDnqCIW1btH8j
PbJFo8EASi7IJ09GGdwVz+E6i7wwDUXLcJgPN2F8ppA9s7xGlH+fPCxSztP1eeidDzdDE6wgFEl3
zBMzTOU1sOpB9xjt7L++YuSTJsgqxWR/4hd4c0EOe9Q7nFt4fKF0hUwJ2yLTPn5fezPG9DMCeE+2
63mO7zctsBFYt49oBXSPH7OjO2EQyAjH3Z5iRNY9LdkSrtnRIBkHPdIJW/wY6ZxoNVwo6EER2OUH
3Qu+FbCLl+ceNZMz6A/ly1YW/Dcj0xNK5uZKGiRWNKhJakUjD4oXs5cZXZ5uSUXWuhb5oMgJlG1M
DKAh9tsCYeyfhvPtvVXQlBrxrGHHvjDzhlMaabOHBfIzBSmoEBef67I5C8ricG5G9RtOtrvlbwPy
ossVgTAsDP5bYpbW0sVa0X0Hd3gkJqUj2wIt0Va202xiwdVilKDN8CtEd3RJPZNdB3cZiFVOExwS
tjYM1jyJwa+f1jYHCOATHPoZsLucO5Z+Ixk0ayvYYtfTwk9Ea717lm07gbdYNygCptXO85TuzXUd
IkdlL+fjdBmzey3j7/3QR+mEuY7qHNBdVaSuOHnB8rm72SZuVKeLsUEzjfkb8z31i8GCaFWAr8aV
9YNtG9HIUo+uMPJhp6aMzd3EHIXF+bRIbEnm2IlZxVLDDGNzBLuXfVocI2j23OqSK1R/IQoPL59d
BAx/eFeaGmGCiF+kZO3QqqzHAUx48y5dMnTlJg8lEimaRdD2kCgnBtcbSr58Uaq+xwxUpoP7NhQS
aj0rN5cS+JO5AdaM/1fM5rEoXJCE+zGLVHWui1sAuXzx2QZ3YlGKVa7rVSBQ5ddSSYnB9FVL+DgW
Q6kehsvgG8vdMhyhCE0nn4p+XitKipprZbug4T2Lv4eCnBT0efGqNW1Po7sIWLd76blETEN2Bp90
NdV2EWXY+DwyU9SngAC/EW0HL8ZAwcMt1/AhyeuRIQmrOAY6ezYdtP8H87hg2DBkovTJ7DO/QQk2
3NS/qFLPE+dehu9XIXfijKRU0nxOJC5PMt8gK1g8ODGU3j6LsEIlskhT2AwsWVDJXqVJAcQKTz//
2Qm1xdpLNdmRtIElykyf6rtQv0UUzokyFKio+33cnXfhZ+CvSfpHgzSWFtBreFoVaGt0qgoHXwcw
MGtMkC2qhRgjdScfriSamUm1oEbMZiKEUWp1gHkQDZodtEAUVppmMCWY7QWR/VGknIzUbH5OupEA
F4nCnkkdRkY0RZGt0etQfrgUaWEB3dZGuJZBl2lYdQO4F00dEOndfWdCoO2xY6rwQ+Im29MkMGD2
QHpl/ndadVbKjBZWCnhSfxNe95a36XCn7Cs742m4U2R8n+JhyU7sNPHeK7nm9fg6vfF5yT87VB7y
g1HgXKKjk4+EDeEXlhF6hrCYCDZHOymyEMAxDyyHl+R6nLJdHZFHKVzFkXlbGeA4U5RpgNJUS7go
g8xqprIf6DCRRe95ElR2ifWmOHDk/xefZE3dHaO+q0nLVOPYuB5xKdmZ7cOnkbZFNPLWz3ZlffAv
k0eZEVToURlnVPsywNC47G+iOHSprGrbIAlpDr7nIOs58+0Jg93r0GkaJ53+Q+MGGArFq3CkQzW/
iOSChCRPJ9uv+xJWXQLWtc6xYc/n21yOEuhVrE2SEMEuaCjVjrekjkFBqcEkgtWfAriyiqn18q1T
yctMNqtqwJXURRP4wY/E0aR07vLRT/iAHvaG1pIZez1wwezGpVgvUxFJ3xKOc3l1eUPAQjV/kcSr
vgnuYdDp/nqQscbyS1wu4gK1WZOud4vn/gWPOSIHyGwWt1/ryymbyuoTmHoNvHQY2JCe1O63AewY
ey4M8M42RZuGEyZQwB1GAU/Vx19VaRxtYTsrdjNHbyVesmFeEnAgvQl8a0gj+/YPa9jwf78DkCNY
b0FNlKqGttOWdVnplLjIh7rw99ETBHlz0tkWKi5976mOBwULJJEZ0qn58JnlPq02sDGHUTPz9E+r
Kd9Vh7kmlFStVpwCHcI+fc5JygyqVvpAvWuGm9Zg8hmNbXuDEAkbGBBz+r7I5xEg/xkCL/FFmtGV
r0K5TdfxpUPaaW3VWfevXw32twfvU1HkmJ2Ei9MlEYHPhY9cmAxcNd3wNqrRJgCcKV2shZ3ElHti
U6BUy2oOY3G9QT1EV+tciH+WMkrcw8a3af+ymCvlB1K25cbRjnWQvbFWbiL9pVGAOX1vgnwFqbyk
vdho80rBZkt1dh5zioHmKzAgYOVDFDQ1eE+7U0p9HmfYB4ZOuCSDaw7dSrDv1ov9lHYpl1QevPcC
NCICtHve2p64iYrOeUA+/CRQzAO4Yx+KI3vtbHzK9z8uNyrkOPgYYNzX9GST6OALBGfpETII91RX
XM7zXkvqvt8nUHKuWgFJZfHJN+P0oq27FXLQ5mrPEwmb+moAAIYK8xI1lSbM7bkR/iXGhjco9vng
hGMCP6YXCNGC++L4TVpVM7oRV0oFCv2Ny/BhNEoKqmqeG47r0UUo5Qqmbl4z6N1v5otc/gXGvbsP
MFnQe4iqFdxwjAaSJ64d2BnFXT/rWF25SUFsjdATi0R0MtcqWeDXhg2EhDxr4qVqfgGzm4CQ+S1y
y+H+UPoL/XvqmboUZF6nmmjqo09phwQZEGwoDcDfPqGxbqjLl+hUfZrQpk0n8Mn2qsITcgMn8ezL
H1w0KF5/bh6kw4dxuNnjVD9w9q/8zwB2qhun/8GOWf4lTa5n4gOZG5J+UMmKaqv5T3aXdF76jwtv
wFywekxyVH6j3bj98A4Q/VPoI9WPngEE+vFcoHeXWA5UXEpTn+Om3juPy6Ac2iDIW4dI7x77TWSH
bd0K/SucV9QmTJW+xKb83GyZEyFUW/B/cp7S10OifSAZbWPdeXJROVsDHW9KnR3J1eyjOEf+HXn+
i0BzJ52LE4+M8AJaXfKvEIw7QDWqh9WzGPOi+hOUouCYSMREGgXXRMn3hHdCt/Y8ihq2eQr5NMIg
U5wyUgMGDhEtkC5yc1iQWieIvZLAhWtlmKlQ8MkVBXkazYfc2zmrI9gKKjJ8pOpCS8aGWh6bl4xQ
fw4cIjDKEUvk645/qsyanwtvtdTSfIPqQ4nWo1D8+/P7ZGTZLkHyR9TW4Y5zsp9gRUm0Znsh/QS5
q9lwS1Mt9win3uueWfknjsHoIvZXrk79xDckcS4d7DZf9NIS/Xu74BSjq/KqYDxzi7AY2iJeTr5i
F88JXq49yFcUfKXIvIR6T+n/mt9vhf76Dhr4BadvdHxNTKeDt/giY9bBYeTKFB9FapTIf3Iko5DB
lsLXM5Fe6ch9pWKZTTNl7UN5tSPm6MG3+S8bo1tL2bNBuL/lzvC3f3TPHjMUd/ZWpfKYCMC2uZRk
gd8K36oqBW/etKTgf58z5Iul+HarrVd4+Hu3l0+9zWJBUwnwbhQoii5RW3qmlOnYoJJdnp2+hJfZ
BbD9EkYDdDnjhAAY3nrI7vFiuyT5vjSX3MDpdYjhXWZ7FozkQAbAXf7NWSxDfngKgcnrpWFgpuZI
r5Z9HD+iuDX7jJBM5rXIqdlW7sYmY+CfmDUSBCBU8cemqls94UxXLPQGgjfZyGyuJbldc+M1p5g6
9FlYu9ByUA8B1K5ZLM2T4IRrtpbSRZnlTo33rXWve0Cq6dhnhFo2IF707MUteKy2fgrpq1sQSwlQ
tyiwOWnMieuRbgQZJWdevXBncmvKTBFJxX5PUaKdxXLqJyYoneaSukNzq1+jmqN95j25KUaGG372
0ckcuYvN6UGD7xJ8O9Ga9A2ZlOKoXHfuSD+YiR8yE4j5HC16vWEpjsLAcAPYybtp0/O3sNXj1gDq
sDYitOQwx+bxWMhQWtmWZFWotkG1nUF4XlmRs6fml4kcqd+Y8rdW4Y7hsS3wM/fpedlGwCs5pxLj
OQ5IkFUlRMdC3oJs2L+53Fc2Q7eMRQ/y5bAE6iuYMCBcLArigRqCLzEyzhqMm6xfti7v3QANziA1
lkSVouIp+nldI19GqL+rL3081QO5hzwbx51qUZpcljStzVLAYpHEMzhQOTPrQeCkiUSA9w0ZWMy+
x6B48iD81iHduruyhr9r4Ii6HbUYgjCFK+CFO+c+6c9LK8uaLMK3TZOccfSou7mDhYRgp6NGIlad
xzAEErTM1WNWdIXntjBaoQxsNwKMqpCK0vUeDJxLBDXE6OZdA2/tBWkzmQqhXzBboDiIFTxnxsLk
9TyR4w1ClyzA9tn89zjE7gi9xXmjCnAUOwE97EUe6w/1gFWUkvGtGdNczX/ZGiHPDNNB8hwY3hzi
l8VzjfgiEuxYUf8PK/ZWfhEhPgiBtJfoHlzWU7xkSCVc2U4Rlo6lm9uOhJiZQNR6PXXX+GUuG35b
Q4f9CoNdnbLz/vfr4gBjTUCoGpGRluRu+mauuCuWutqT/6PkiHimWrBoqttnJKjKKqK8xMTt5Gku
RtFcdHMF4J2boIU8e/rFn808LnP0ZLMrlNsmzhOnGACf+h2PlmuK61L0CIrcQlWAllR0xj6slLEp
rV5x68lQMoW48YEXRMOs+6pSohv5YQADHvT1IoDnpc2SV36EKncf/XYwJbDd03X7+6iAN3pBriHq
bczPYJgGdXMmUW9xbveCvpjspO9lw/F/B3gfTEWAVhxuHjon/yno8Ck6JDoYeIL9JuMbaPkAHHbN
/oGtLNyhFxHLPlRzBw5HthH0d6jtEQNCEy15BozcjPEpNMwdsV8ma1di9aedVPuMaX6tGGwjGC+s
zhK3ITh+uFdhiE//VB0R1uwjUkWmYlT0OgRynmOY0FfG0TJDccCMQvE/TYJFrLPIegxbz3f47XQb
vItLIzbTWPmmo9YukGfwQqvl6nZFn++hEtE5C6DCkPL05rnJaioOhN2L8ZEaQrr3+ZH3fw4a8aLe
rtxE9lzBg9nso72aHkO79qvSH/FkQabQaXBA/7FyzxhQ3e+kgrbp/jWQ8vbPQcxiWgcEGQuCVhpS
DucNb6eVn3ThzkomBYvOEX2xzJ+r5EChqqYpOC8rddaSoaDgcLq08KAUCsrGi5QBKtIgl4CDh6xW
44iOz/yLHLUzK6REOZ40bFZUlCM9fow4IMXOjbDmtznStXPKmPSAv6CucP31yh4vxZWWVMSsc911
Ud325U+rnQuFYJCxNAc0BkxGMaT+jnU2/lnmzomPC+ISDf/QiPxjiVYQ+ccffN5O6jJqSp1+6hvB
5gja//gHy/cvFjkEaH9pmf3vqrT7RNK+5iVE7EtSckI6mlWGdYmc5UvT3isPV6Rue9HE7dbLzUA7
W1UEES2Lxea7TGNVESSQADUJJc1wCSWtHfgbYjod0pWO2w0ZXlao0xK0SvAe52dECrG2Ad+Myg1o
5Up4dvh6ZIOdRQju08KuzhvJsWq5a5ic++vUZZtAsMGP1/2WHryicacYbRyKB7ljrC7swsxajhDF
uIidPBlWjwrSWEcDBok75AswyHyBGeDKw8mpJ7n+T7Xik+E3nYNQC8/NsX+W4PwEyHp1RfX6uI6S
OessDQPUAqnKNHdqV8PBImizx41i2jPmW8H5GnuJ4pbJcEtPkIRONykgKEnerubqtmQNMFP8Qnc8
WAGEcT5riPpQsyJM8a4LZ0BZYYfBByW2z8l87evBIwjj1TKtR8XI6Lt9VIogANvx7l9q5w1GA9Bx
XaSqPWm8if0pDyK9yeJicT6xWs6dEQ1oSbrkDJgsowOchl6f9InIW2gYDr7VvSkyJT7R/mTULjBn
UVBKuElQQ1/LTEtTF7QHFp8MY6nPhJXYsKgXEXsnU2rUaTal75PzI1dVPJc3ncV5NUC0usQUfv7a
Xu7EnhTZu7Py0sAIBHJaiEWlmOfBQ1I5R7/B2nyP9HUntwto+xKLue3Crurp9snJQAk/bPDYyU3E
KRJVs+r8pc5CkCPhjRZgO2NJmBaK9WwFr3N7k6mafZf9tr/bMCAxmc7ER2calbrs4ge6x4klHQFE
cI6JZgsVyw4EZ6DvB+8DtmKFZHn+SGfXB7b3iZLf6T2G+SQQYfYoai1kYNGFdCQ2P9vTqyAHpNdu
bvBiLVGiNEKVvVlvXNZ4IBCww3i24vTEHp5+1w3AASo54jkk71jHjifdR6C0Tqovaj4yS+OwhD/B
f6ZATg6Z0moCcd/zw9yaWEmlpNc7CG+rmtvfHW6llJbzmXjA0pjT9j8PYx8+GYKHFVSPWBsVxEUK
CENYk8okIcfjvbcliQl7fyWFjVVRE+eBgfzefKnZEV9a2eAtNlI3JrOGmaEIUmrCbJNqPJ6pD+PX
l7CKIYzF2wwCRRNnfCMXVEQPqXWTjd3o3LsRpobHVLU7JFSSxqoQB+1kzT8bUpAdyBGX6IhHdSOg
/R77TDILIepYcEC8+UM3gSrGbLHWaXsTxX0ZMUWSqjDEsXV7Xrrat3eO6QiMfK8vf9LhWszAKm7t
BZsBOYuuFycGz5UEnyh6bVx7eUed5vpy+kx4aTFsb6KUiE1cqDWX3PaUlH1FqoTBFeQTABMHz8yY
Nk4iBJV9K3ih/zA1CvjfDjke1osgoM/0wHa9yJXtROTd245u25u4yDd9VwxxEN+LxKDmDtn1hwVv
Tn6KK6UuFhRAKHGtnpEh1cc34J+PD/T3JSHVI2QcpNVgY2dTqqlExABEQOhskdky7fTZ2MNOSY5k
I9/jOgE6cRqNclLtrVVxYH69VvHFkigN42dVsZ2DzIb9e4EtkGxkzBQ0h1thaXR58/kvk/JEeA9p
wQoAa5DPICNIc+P0pMxFZ/P+/NnlAuootdiIro8PTKf6wibEFkbR/nVjbQ9aqRqF/NmNtFTUK/fo
d1Oa0LQJGkOBjumxLbL7OSLX9LVNLsFLcHCwu/DmElinisoWg9cyzKzbX1suHPhy31YjaOgVIKp7
ZisO2PPkB3eNgHaeuTW46Y8T6ftRm5WMvu8IJZq8od504KIxMoDdx7zbLy1vWy9lnmKM1clsPJrq
gLvEPDJCC2tNSO6lTdBNxkY2XLRDPxhP0sn6oY15VBOoWRLjIRyQKkMkFYXp8RbINk3IRR0XVByL
tZ8cNKsEZhSnl+G7jChm9AYhSxLUJNRxtE1zCRh+gamKphV7w/xUuJ+wN1682KZ+iLR3txUKohBE
ZGyJa7FK17/3/VaF39lj/FStT+6Z3Jevf3jdXp/u/8aS19Pa1yKUOvMPckMcYlCvtWClHKqtbLAT
JdnjglmvR3dnfQD0F4wZYAA4m7UFnNNVKlf5UTJQlbE4dEsjV/kNf/tjfXjRt2f/HOGntTb2rV8Y
0qLlTABx8kqDL3+3OZgoBZ/72tSFr+7itKlirrDHYlZ5vHJOsKKWJILOPFkgLf+5U8Vj1p+ihL3c
KX5YlFMTTjhNUr8Q6a2usHD/tz28Qxb7tm9GoFL1GAobD08y95UlDaZhuq4LtV1HjxpV6MDZ2dN4
jk3gtXSH4MBohNuWbkpogLBxuBI2Sayq1ns1wJqhSYihRDJNmPmweeMkWtZnTmOBIQygZdyKTXX3
iIxfHKLSNVcVwhfhGTxSsobT55RxJFGVUkGCVZEAhAcbn+DKK/BiXp/Zox5fHEV7HV4efjrnXyuQ
jtWgrSwopUTOQdrAaPZehhxg22t2LNzUkr1Wqq/UOnNifl+HznWzHu7vhrPmyZKUZNykm1vWI1x5
GQVAgEmdNVYhwrsbewbr/JA3pAY/I4wdm+ab6Ec+urdJauEZW5IaYK74HsP7SgBX3FA/RC2cqX/R
ic7KSRLxz5tLdj58a6WP5HvgsFluYPOvq2yC9e3EPumzwe6GPixIFpGj2X7RWbi6CnzKTL+qN3kN
1qMkHvBOGUl6LhViYblFTXrZsKmkD8VcGrZAfdhSJdIgebfjWPmDYYLfH+8jttcu8IMvvXnkne4H
YIDMPL/dYedIDR17qsc/cuKBfQx8/tJWcwkzDcIr1MUtgqOMkLftWqJ5MmXZEiSCub7/1BHpDBdp
cSmBm2qCK10xpE1fZq510BAjipAVZ6OKZk8bLsp7C5sv5PFh2puSJ+X8xmtA2ReMAiHmRMz7plq9
EU5EjwJlMAoegnbtEJxCXgbs7CpHD3jUvfmwsrq0gPPv36dszsESyeZxjOcK7j7b/DFYjsnsfUbK
rEAHDnwxidCI7yjxVuTKeKhiACyMHlYveaKr5YpQlzvjLB685wWlYV6Q4419adRZ3mdetPf4J5uE
JM9EMeU+Vi5Az/Dml5qAZ8hDsq+Rg9wfvzV+rJ872dHjWWFi6PEq4IcAFis2RITZLRQyQBcVvttR
j97gQ/toHQu8TwHvHwxWebehXi+wc2cCu7DxnFaPc59ubYvX/kf6uS40dd35sB/YvoecRtnZUc39
iKgt5Y+OBqcMzlEIP5WG6tY2GWcC9VURrRc463i+F+R4ROCpoyoxYlfICBNce8KSMJks0Gv4wECs
gWcLn77L5Svc58micalx4Z9Kb15hqvs+/buuOTSbdha6AfFolqro3JoXh646B4XXuS0RLGipX1dE
ZyegJ/nBHwZTdkl8V2NjcSEUL141RF2Xm3ml6VM8HW5FFSXGU5o578xICnGPyhMz4LQZDLXI8nRB
dSAZBct4PFkM4jUlpfIh8/QFmfiU/QLBbQJhFGXHpOkZ0f/XLbybfBOLtI3XDhS6+2B4J0jaIHmB
/O4BgZBumZjVYEJurJw4OiK0xmb5jpsMt67H9KBG19drNM937BirmcerUJkQc34ZHOVw/CgGWviq
gFebc/reWbS5q/icyizwrgeWy/Z93wSoBS3LLXu/e/4xT0G2P2MCoyUlfrO5FYndovp3MMM/E4jc
Ti285y+rFxRl+Yw/sqhL8nvn3cqz2ecUNHLLiGtgpOWZsenLwl1dibt+mqazhSIRoCbCCcdYJjHp
2lXQmUyHlqnjTvLyLo/DtchYxbUFKLwf56ZF30X4+qOlrX5rGDcSM2SjiAI88jzhCf4uAJKM/v7z
82525ha/lZT57OUDmM3eYIp5ZknqSX4vRc7ipa/Tjn4xbeloaDz4oDF1XpUNpALbUKnNBNVwzLLN
CT024DrbMwQR/h/I0vZCJGU7Qg9VX3lKlbf9U4XRExPKLy6bYAKxstp1pePgM3OxRBLD18xz5h0Z
FdbmUUzq4TbvCOAel6oNid/guNHkZP6RV0gqmDiseYMv6xA6kUOalAqEphUMaqhouuGxTWrOEe67
f1DR61pDbmztLKMU27wFavHrnV+BZipxDKFi3EJcWDICBn3nXMc/n7LV1WDrAtpLt7QsYGP2Si9s
kI9dcbm1GqKdqRkf3u6GNol9XMajPJDHpkTJolIw6MD47Y2xUQc2pTbaLMzK57NS3myhmr1QFskv
5KrySvmrC2kU++n+c/1ssg14ObOf7Q6IlQ/paiHPs4dGWjhj0iaBgKhy15EdVeS6xpSjt3KVUYhw
IeTaeBCVHC9JiYZDxrrND5iaQuQcyo0C0jJfoukc0nOTH9DyulbIsFwIBDt8wX1jF8PrCYeQcbJ0
4uqUlPt5/luHeIkejQOV6B8ESyv/T7N57EAKJIkMcAJV+B6i/YoLPDIquTZsTv56/kr9wHyTUY6f
RQH//wtRhI/fv9ZXPFH24Qqj1oUTeknDi5f/rJKvVegWkKkQCuImLHXzMxiO2YRIyom9F0upEhZD
cASUE++MWTqyXklaHSp2PkmDvKuTJ6Y6tO+qv2/J4GxA296HT/uIevrgAVhHK2MTKcWsrdm8sydA
l9jeaQ6+BtbW7lfoR4Xto68H8jaPfBVoa3jokiJXe1GXqSJ5yeUIkF4vjoIL88Jmz1WJvksohzR5
1vnuH7GGsNA70LP/44e/kWoNzxyoILOlq/eJ/JRgMVhTcTfo1MRb9Ak5UPn0nImfJ4Ii9vyWmqrW
kE1CtrS591Ejo37GbvuAsv46DoTUYPXpoceVHi2n3x/4LC6MjZ+C8ZCtIKR+ozpyyVJ0iKVb6O2K
m1MubtRLVTnSfZOCgFZ7ue9Lz3uth3A8NpkVmOEjy7u7bRmGN159omidrDjhHxCf1xtKUkM43BKE
2z73DTr59tbolc70CxbjXMf6sSCDGz1+ugNKsFv7A4F+2xLBIGAKcHBWGF/setNGmsEqqKLFuNsQ
QQT5pljRm60jBWNliSfCYSpGgqQ41FASVzbMHFQ+elwmQfdH5ah9ZPWWuo/O4cn8acaNDxmC1hZR
2eD/urp7TuBSgRLEhLOTzrPgHNWzZBdtQ+QL3RXztVJSxBqRgggYd+0JIyHD7bvMSQSi050v3riK
SgjdCF1YhXKLuPDlyN/WRlyqZhLxOLsZv4QDf1uvpn82R/qmkwxlsA1RzkRFigPbBDgnTGZLR2Uk
2clX85GaW5lIb7tJafAdKGK4iBBjHsb/0zXTpBds7hjKUqmJzhr4gwJd/SLRKtIXNV1UHEkza+f6
rjDVV4uDAabH3UIF7lY5muLLmTeXAqFTSgIUt77TDqjMu12WL4gnnV11wVsIm0V9n2pBrvfxPq7A
Vnhj7NbVOJo6m6sFKZyMvC3EKdMSHAf+tDF9hGopaMfWH9rdY/t8Lcn83MKoPjVYLE2R92xzaQ7P
8c26iDsIdHoQZWRHuVsbkxzEaRyVIE/ZZBjmyeetPqANsNpqR0YUjBhdz3rMld0yhFEjwOcHBN/n
vur3fBBaFnsRgzXmED34G54cSSJqHqp9ysRJ960a63pRRFoGVcjiTUxRZvBURaHiw2L5x9IH3TCO
ZBn+XO8ZoArcERg9Ruc1X5zh9zn+/znZT8nkWsF+KLe1EkeMPZLDBIlRVk9BqqpQ6YHYo1SMKlvp
VjCVyxVrmO1HbpJF2KzvPG6litq+mh77w6YwckUPK4MQh4EQWpH3ULETDLms2M8RFS6UGKRgWGfn
EVMDFJlKG0JkSSpEhuW0Ak8txEZoUnwmpelmHlHnWc8NxszlaMqyoupLfUurcGiA0+oR7q4kLGsq
FXkE/eeIGavUYZgNiHgCIGTpXN8fW+BvjkXyo+IAdxVZfmUovHUjUDoKZSixBgJbkrYNgr7yNs/M
3S2hvx7Xxy9QstPNnC8gpW8NPcZ4BHUhmJSiIHgHLwr3ncpXJqJ+Q0y2ePj2DKgSyAY0+XrawAZk
oOy07ZLHsseEELUdvHHGvy9EuCmDn0tpfnR+trhN8AtE7qMZzHPhpCnNI3OFxp5R6KLhRK5I4bUM
C8tAw5+o654lNss7lVtyaD9cuJrr3yy3H76Q+doJZFW7LuFbJ25y0kdT2Uq3bK/afDNE7F89F2WL
wDdlmv7/lxIi5bvY/UktQTUggBiLM96+cy/PmwPwNVS3bZqfA7rpvgclayWbXLsyzYmNg8FFvIvu
mAoTHSqz+JMpGa0YeaFZs0XFuDIF+z60OvtSY/u4X08rVlStQrDf5tzOnCezqQBKw5Jr2UAxq4Fd
OOkLewrEbWDsTjZqaqkvym/LwT/UEP2GzcGfJp4HkPaOGLEKzJEkV2Q+tgfq58siDOxW2D3D8ijl
cnvYc/pk0oweU8smG4+EeK5nUF9CotUnchnXagUambheu4bcRvBUJxTY6rioufW0z5R4/dZS2OJK
0C3s+6xRk51HHITCzTE75yDZ6ScNBXCs/J9XKxGuF+HZTSSGpCcjUvdtCW4Eo31oILFtH7w8mld1
IowPx5nIeSwADTL+ZoVPYKJZoYhm1Y3KViNZ43gMyWm+E1GuvYeQnABXwPz59eaUd4/0i/WdLtWX
iItvCfDwqLYJPEkR4h0fruiboIbILb17/z5G0Ia5Rk1JYcUoEwdd0QyVK1EJTagRZNpdP+xbXepk
YaiLkharMKWWK1Lxxm7N8O3A+K3DbpTMuRNtjUqoj8oOscIZ3l32vMxX7nEDQbxlvR/ZKMQwYShQ
I72XSrYw5OBORGiyWaLUzzNpCfi0AwoBv9pKEqyk/ejhRFQpb2FrHCHVKgI1FvvCNOwv7SnnBjgR
76UeCEHuX822FGVouY486uzP/5WaW/TF9J7WwR4qL27u282jp7jINA2SDBH6xul4L3C2C2Ird1Rw
nIqQ2epj4uwBOE3PxWA5H2m0dUn55dxiXIuETPs0n1b1yvE63To5Xrn5bOOVqhyKJDPGXFTt5QGn
BJ+odNGwVn/8rOcq8jTw2xYvPdXrejpJQw7V9haSwuYUzV4dtNR5zFO6qev7lJq7TMXdQoxsU830
G4+ob9zEzS11aG8Ts38879tidsuOgOnPDzRR7DI/XvRR0nGez9Amg+O/dQBuDcAPmfl7WYfR+GSJ
8HV9IKc97YctuPUiaLl26kgZBx5kNTi/UEq4bScmvI6zR9SWAokRPgCkrt3toeHfGY8iE3/YNsNF
Y/9hVd7JXzLLU6Z0pYuzWSKoD/FA0MwgNN8wn/wH5Zx8Yeh1ErnLFMARKEmdsdLFZQ8vDdktns/G
V8aRaGCBMkt/NBnNJ1SFG61aB42vijX0I26XIbjoIj6TM/hlP8MJ+W4yjUuttSUBlvM1erDZ3nLM
WYbdZKNiDwrO6IdTowaxMe2CpyfqMzezzxU1h6RdbcDko58Z25HQcQ8z8BmUn/rE0O1mbpScQ+A9
gJpeSv07NUhNdle/jujrViFbIYkydC0wFOzblBzkNNh7ZIRQtUCSQYtLNcGjtxMqDBMgDES40+t9
qQk0JRqqhG1v7XXia6oaEDZdsxntptcRi1iOV3CPRcWw4HwIB/kKjagDRiXQh5tzL400kTUsnd/2
3eEj8vT4ctUcFTczgQK2CbE0CAHafyts6T94bdMO6yPVi2u3YfA5EIfip+V50HaEDO0WQGZRRE4Y
hvCbz0pTxpMQx0OIXC4T0yjPpgxrL7rhgut/rhX/CPC+bKjNc6OoSPijjxGfJOfN3PvsuS/QG5Ra
biT6bnEMa40zf46Jbf72tCYh4kvZA7aApXySEyWzaRi2QOLKlMTMDBxCOaEc85dZTQrqCUQmpLRL
tk8mU8mDYFJ3GUvMGibzghao2+dGxANVIJzY+xL7djOTgNNNj/aXkxqgvu/QybkYTDdyYUdhm4JE
13Iq5OINqCTjMLuznVVk0MMbTw91QU/K85rjMEUK29sb+AFPowtmza3zNpwDuqnDDKHzsO9md0QR
ajdJiLW2xlcayyl7KZKeuYagAJnvm3UfdKdzy5Vw3RCjm/GUHRsl5MnpbYl/wY8qk6Qt5+8eYfWK
2FvPAriOLixVQKEHyamecCdbI2gno9bu7InxunophLsEGTotqiPxOkPaNDdtd15oWDcwPYzidaDR
F7UIkn0KE+2KksBnZIxsfbm3R/Z9HjGLzoDy6hq2cnl8Y9WkICjdfPf6aywORZQhWABh1jF+Nw5e
Yd9X+Qx1EA3ptpOLmISFX3s2wDGl2MiSw/VzQCRIUd4EXjp4hxp/o4JPOx7bJ3VkO321W1TAmhry
2WKO5iKOqnAqkkuedCAqBXtA6chC8YQqGOyvfcuwJDWIAXniSmLX8JFOm5Ix3DKyE0tcLLJSeSFA
oP6id398W6vtkkNqV80nb3C7emqVsPgndNuUq1GgwT54e/2Sw2o4e8PliO3Cf7Sc4Mn+xT9OksU1
gdk6GQkDxmg2Pq9cNRiet8fP36DQqnBxXe6EBTF+Ijn9GWCf05QjcWvJZS2lTP/yTgPerH0K9Saq
3AE5OBG0KRPXW5kw7HUotrE7Uhzsma33CuzRaK8lDRbM/pnIm0nrkEwyMMzKlQ+sbJImxHBLOVui
EiqCJoanCoMUbQrG0RLxfJVUDm6wsXLPHzVxkJ4kvR4JsJjjlqwOjkQh5P6G5HhoJd4Y4rOZxvv7
oLNwzltQe4jJRxdRZkGQ1H8AWn1+kGISfL3jpGt9Li9B0lfh+vVlbkHBRPpWuYERugjOjfK+TZDi
zaVCoyuhXibn2nf27illvgrdYKBJ4WOEKzcwKNGEBOjfq6TMXRnZNlrt9ZFmNUiKtv0mBaOdtTwj
3ac+4yGxvzSoEXyhDfRYV9KcaMzWNZ3dNjOFMZDkaYnqru6NGOKD81o06LJqCbzcSsu1p6EBbO6o
lMd9XtyUD4d/aKkalCGaVz9E3V6ub8bpr7mSp29D8+Vw6DaTctzM6/TktkwtPGgXjOW5JFt0lfzo
use6p0BANNHgyaNaTvA2gD0vLko41TC9UxC+OW8wBnsG4hPs8ZTf8QjsOrfNFEBQ4Y0S1AdZztT4
paFMwxNcSwbgabXjQ0N66tZQ0iaOyK64KPkD9e1UrgVIcbgKHIS/4ooYQ+2eo8aGhzEQ/xqM8pBD
9DyS2qMVfAVXqpW2kWGhUXmfXjw9/CksH9LCzBNeELV+0DEgTPy/m0uZXZIrPm9FZcWw/BMxVMGo
tHabMFRbSp1YW34Z1tlOzS95uUTkufxY6lzFFfQwRcHca1yKFC0uwoU+J4+KrUqhd6fGkOUIwENi
lbCoeXJVwPf09NcPImDZJMbOKEaIkLymX5mbRZl/GFTNRIXCmNkjeQdwUTMyxm3HhUYMKgO9OtAz
SKqCnWpKw1i79Ttex4Ht7U0etIgYgXqRSyRcVTwQyw4JcXwMMYkUPFB4mKN9OyizhsQYMfEYnRAK
h6MNZMNaW7gMy8m4rdrazvknF6I85KMW1KLQfkMRoETLlWf+on+kM9/noQwlXUPBGVArE8fDyeXK
z1SbWBfeaqntFzvePF16OgAayhiCYFY+a5MVQL/kkAoRNCrzsR5kXB/gllA0pKbDeXweo91OeLc8
xfnfm0JdAzU8mHwuuA3+WqF5wTPFG0w+YKnsEPePcbiEvFWSELKKTcjPh9oseviR6J20vx5HOkK2
YH/u85n0OSyRq0AHjHU+EyZaFAMlAqmiYBq2YF334YknsFsfo77cjDbJrDO5c8RwgvhYjWds4oLy
I4fL76RG6mHJF1uU7XzzfNRdacqy/w36wKhBOWDPvJ3pyf+h8JG84zUGt9xzgo5iZj/UJzKcqcNN
Lnb343FXm5IDIcbJYi68wPGVQ8EK9IA+IjGjoL8xDyKUMi8+OdDBeDKxQBC0NiSq+7IAKrui4keP
qSp1sOKZE9THbssJEpVMOp64Xb99ZJ35WwpFUaJSb1SflUx8HFso6TLJoSOxMjPs+043QopZKwpe
gl0kUV6ZgGw9q/dWsZ04doYqmsT+9n2Mxtpr0cR3A+6RtrTk1DeFU4viJYiA3KQXYzrc2uJbOVZs
HyGnFkRJlV3S4RVPDdmpslwIkX+liXCao6gvSHpm6YptSYZx9Ru6Bqza6+Xwoc0ut3Bug7pd7M8/
bvW8UmS1dgjTyYKxATNSjxVThTiPd4QILhSpzNJnJjzXw3NIygK66OseAvTm6FqAtnrMwBODAjE3
T6kfVRRgLU9QYRa1/Wa3XoQijRIMBb0Sy14aOhDJfEYXTYu/gS6oGhbHBA/MM9+oq3KNVRTvoUcC
NcmEMUD2vm+VmcUUmV7fFAtL4IXzQyI0d1JGzV2UEaS4HYeDESBMd6oE9Nmt4V/XIFXpdUP+js9X
H29hLF2P9Nr87WvkXMtsc3H/7wjuViD3joP5wVMfekiz/OAZwMNSJV6cEwQLtQLCPz9UGCHiTLoU
LMnIvoe8pIZlzvRihqmsuTAlgxu957aOFW0qsqa0OKdkSpau8q5aiAB4sQAhd+ZipPvLrcqgyFEe
8cPFdDRMmPqaZ6Pz7AX9cULRBrLUXJQrYJ97MmOzvhuWmxuOEHAK60cDgnljnlb582LSqvOfdxSI
cJONdTbsx8tida9lu2Ga1Ywu+aEeG73pe8xXDno4NHtsnNXoiuxzgemT/55O4ZsC32iLjdFR3Q+m
VEFNqxVlZdVe4AXUHm5HxHaPDd+mqAQeFxCvmTCiDc7YInxQ4FiCR5jX3EnfXegElwDryRMNK05P
1qEaaCwvkfHmX3VPVlNKuLCxVsLx4Hn+cNZWTIy4D/Fzque5BVGl5r+/1G3Yiwwp+Y+WpuXX+f71
8z6cQ08+9lv9bUSOX16HKDO912V2Zx32EJj50X5YAzNvpsWs8LPbLdE7+MGAt0208tYT4Lss9pxt
R5ife5L00mEXgBHmm3oOdGPJuGg4KRiDADt7ektOvCEaU5uCjObLFGXYdiOAAWPJ6izrFF+3gbMc
gLd8NxCDQv5hDAwv4CL/cjwqK5U5MW18Doi/A4ipToETQMTbNafg4wIQ6Dz3utR7sqTpQI2bCJp3
VeewN1HKLay9fCbRHk2vG8gQMqgIxgh05sn94MV7tO9ygIP6ZwT9v1UZWNoIdL4YKheLBJ8pC67T
aF1OLpOSP6uMJLYn9y5jiAeJ7U3A5LQixU27ZxI704CaxqLg1BbmiQW7SjtrmpeHNQnE3Ls5Z/fa
j08Q66xD4tyLfCLxK+TlxigmUeRwTd0GKqr3B2Aj0YIctNBzEHwoiYgYCJRG0N1G3OvYF9qUVZaZ
W4+4Bbw5wIoEKFcPypogKVvuU0dcmhlwrtMaZELj6Fe3nG+fITyW/qS6DxJwOtBRpMgXsevuKonb
qAdlgAePWR5rdR/AK5sjxJfRrJvRbhsryT/xWVu3GM7izjwjhB4eJfo7GqufJU3NLi4+fJuA2DSR
0Fx4NBgs5DlkKOo9m7X5wv2jgLGjTN05pung4u2VzlYHQlKsG7R2uqwUhldij8wxwKkSqX/gwjpQ
haFGB9Ul0YCo7IfgUA3z59bftP91smLDg4C586UYUvK4L5Da2izy4uQ+xS2UraFyVaCVmQMjFQoI
d1Tg2aM6YBVb9JaMkq/ovRfxRnRQKDIO41jqIXnY2LEQsKPJXMXRVzSRKteFTzDzMlHwl0NwSgkP
qirnQjPLlAw4eYlGhh63kN1zueVxJJuISRSTtv/j4gpFTvY9BuycMmp9sxhkywHkrT7rLOIGiRIi
E5leEQLGopGuFODVV5uo8IU4wEpYYN57JmU80VT7OzycDshzEwK3mJzESIP03kKUD8Bjyz/Vwx7f
+sXgz51mZgNcK81juEbWKeSYimJdUKsURDgPCKTgMBOELFwrL33Tpkyr17jedql/PeAewzlMrSBu
4CWqDZnLbgnM/n2fzVRPSpW88/rrnitxAPPjBsG+XIQmT0phfCxbH15WABklhLRMySeGT1iJEbVz
HfyV4Xoe0K2r8wMn/qaGtXepeGa/kA5CNYUFPacPC77FbxoUzTcYg2cBKsYkT8ldNjmfAxhEAOcW
vm9vNot8nUMmo1QMj6p+IDt+4N3kFQhcOHnzvm1E4PKUvvl1WGZS0cBek+gih2VwniZDcwOpcJgN
p9f9ZCVOrgpNxBCbkHaQ+gxQRE7g1qgas/Yo7yEyFfeFJMyH8vTnzotKHfn/QkUczlut3k+jSmS1
SZVziXck4Dy0sxg6dLYt8oVceA6XZgGg3uhdcq3/fCZLHl38if8rM7mSzSlDB47+NbxBHig5KqJN
HKf9VaA32kPNALzf6Iqm2NjNdJyHps52DuXPSvbS3i+F/RGrSkHwi2Q/ejkA8U1o0qyUbdbbS2c2
vFn1QTGAkjS1RgQIJFOSrL5N5pztdicH9oiXBuxJmRPeQDPAfsHBhhPdfaRZ+UQuy1zB41o356Ao
q97ZYrMXOBitFj2/HtUE6WPNvVaR9YOe8UABirFoCGUVYbQPB/M8ObGQIKoK2C3842SNnaHiTiyn
GJzv7VOchGmAkAcW84Ernyl+MGs5jg/zAh/ORX31N9Rei8C1CVicMiDhMMU8QHn/vUlWFTAtsRy2
jG884d8wvR4ZNsFBDmWBeQ8qo5aPh2ms/FDo07Rd5GJQ/Zvy7cMBAxmZAL40tkMI3apRQXaVaexY
3uY72Bxnz9TgXwpkylMNi/2NsixA+72Z0ubFe5xGmmiq0D9r76gpYeknFM+h6QKarzEMb2l7zAif
Cu3ro4CvjxRfe1uiuJhaGewmx1d5ErOBiN1wvCztbH7mc0mcF6ZfYiUwxlpYhx9UzYze/XQKwP/X
/qQdNm9QFYKojCh4M5GopRAgUiph/Dv2c4hkRYB+sDmVSp/n1gmON3Z+qTSXSVhYlfmUG0JOSsOi
ad7bFYFRH+0SSgoHMIR4IaWBPv6ldU60GZL5UrGZH4IW4QIJ4WxDSqzhE1tfSdsK/xh4z2S7IciY
aatiSUHLSWuhTRDys9Cv/focmZRojuO4aUsEvtCUfXrnf3rcIwK7h7khmiMa29oGJnamMuxJdSvs
4Vs57RSuc96It+WCljmmBNB3ndL48wSFPbyDLz1esd5bjd7sZiXFb1MJK83O8b7XkgGCmBRUdhij
JpUsfbYtv+EQV4P2hagw8YqVJhNtWS1aUPCY2vWZjUEBPinHuTT+WpWg9I7+Ix6NKHYX9ouKK21m
8nScJTX66ToCudspDqbZzJmmlODmK2J4r0nsaaBovHirrWjKsXSyvVm8cVrziuhQJ6jUwgFQEDrb
/jmdnCKyyI4V4Z4EsVFV3PVI9/5tYNrinVHe/67RAx0L07r63UGgTIwoKBRnbMnxswr0Qt3t7boF
5GfqwtaFDjZA3IxrGuNSfvbJ6khivlwh32hjJhOTACzwwf0Z/WaDyQpvUceWgRRPh/snEG5MPI7r
Fc+HGEJUT3ry4iYrLoekINvF3BYgUVPBpfEHMENeZITgUVsLazk7IkX+huTiktBGxynQ2O+nFxea
g+m2lFOzHT6TQQI3k25KsyTowf05bikt2eFH3jIPLLr9AzTH6LdFuY1olILbsU0OXX9z1pwrJRVq
Yc1+EfLme5zR+ArIs87e9ksIWhb0HwPEzmAy4G1i2mUeRrP2BD10Ve/4zA/GEUeNjGSwqJHFZKpZ
1Jq82IWamRPW9AuBjjXmJ/EwzLzB/cNa8FnOt4fiwrr8wQun04IUemDeExrv6RzoHiFkB863dflb
bgyUC0FZFJuKcMG2+GNXWOBR2tBJMIPoDsrcZDLyPsSTCedDCCfDQuoebd+k9Xg9Yu7BUFdJrnme
qo3fOT9bXnfOVJcAIz+ZuND+FGH+PRn2GNBWjsfljnY4nbO8TM3KgLm0DFH+KMmzl5hC++39ponw
EiLRS0Iv0fhAqEA/gRPJdBwJ2iFhMe/kWy6hTYeyEBMxC0FtbRcAlUghNwnL0SLjjFfWjUoAJlpd
4tA2BkoEaHUgiclU5YEUxTaEWBqbqEKuOX2z215rYxgBIe3G9ASybyQyAnLR7btoj/XhZFCwg8Ih
DvY0NQmEHI8exNFN2igDQaLkKamNgxZaUVxmSZkfkjCmUEDbTxmutSnfI5UlDdjhQDri92Y4EMYQ
q2dw84VQITKTAQ7uvK4Udtyw9snA5XOk1TlpJcP/I8JnCqGji6WC2ZwpZPYvoXX8QT6/0u6VzNUo
UGWPYioI9Jl4r6lCJDZghl3XrsofijzvBu/2fEYiu/u4yG9j3OYq5xnxekqA4S0mFVBMV95qEETN
MiCk7WHASe5pFzwTEFAtNkqA1tENsa9aLk5CXsDc5wPchbbRB7auuDxayxznEAgrhHVXvn62pU8Z
hQ959FUt1+2zNPZUoG8fHDc25HSk/GGZfzYxQKGc8aCM4jUsX+6VHKKl6SPDt0KjuokGu/lnjmZX
MEubxFlDkaDr9m0UsbjiqWmTQTqp7i0BymzusVve2WNJ7reQraV5+qB1GQ7r4mmht0QORxpcaxRm
zZN2MkHn0gxXI/qE2VpzALEmR2ymUMcbvuDIYlUMlK9Fmmg20JhP5fd0rbiV77FgWNxNmdPQwJ1w
HGAcGFZSF1PKt5jVjkIFy0bT9x/5K6V4WZZQPglCDyJ8TtlC9Qi7VTKEQvd3jxf6P8/aifMcop8e
U1Q9/g49OoWBhpCjtcRIVjlSSdFnWzFCugBAh998cI1xqto2SfwRyOdLQwrtYH3KnTHYBhdq5xFd
V1h/u3JAGSsyMyvpJRAWRdTxKqAq8+2jEyqM6NuFOhJC/ft/O5hMbo8FeeGIe8fS2n+aRvjJsO2H
2NZumbuD5KlzWFz+AUIV13QB2ZtBkJyHlsy+yAynNV9VZMxkIDTBjMAjGK7viBXzM3UqYEDNxB2Y
/zVz4k3UhX9zbsc1R1/VKwQGDqwdpOzWxWdNHCaMT/Z2pAbs1VDEIvPAMvCKQeE8iZtKkr4TXJP1
CEA/40NnjStcWdN7QC/huKyyLQNhNDZcXBLptCfPgJcb6dLiBxRL/H9MnTDB68/l7RsHVC9FTFEi
Q4sm3aUPHR47XuMrRuFkY7bnjqpN4Uc0T2g6sMkRXKd3dezbaGVAs2My78Bjt4ZZe+0f4U/vL7Yu
1oL86GryqsTe1qywOynMF8ESdQ4y2ZgVTPelbJEx+oRJIxcoJyRju8LeIF7uGxv5KkBxIszZQ+Jr
n+B9BtyVmM4G8SPLIKHl/tI5Yv42DZbinRugQmsFbVLOK6Ltfdqes0TuGYFQTzkrtUGe66lsqnEM
3xfllLmQPf3mmYvy7B0mvCAzZPHAFaWdqKhp95qK6FJruBxuMiNOxw7u3PdRI4iCWBX2Tcrr+0/g
5W3xIETLbEw0QIc26sJCP8IhntdETRutVrIIIJLftPEuxYrjRZZBP/1MjDr0+xPWqo70aIF2L2Ky
E8w1/JhQeZom5aApjMeVLT8y21yhDA7MgokR6ApH8BRzTVDQ31VpL57CY2JmXN6AaXgAreFa/uLd
rNoU8bAGNS6TB6AeWeE2IyKCHWwdBfCmt0j3kReB9OQPoNat8QB6UE2eg9xEmHyWEMUpf2eFlRlF
7Z/VZ6ruyD+H7DyJ0hhikj3Xax7ExgHhPynCB/QeE1gIdMcyQBhw2tVo89vxqiS/W6/5CaV5pzs6
2kzwe8aY56jzSin9fLvFXw9yG8Yg7belQ9scoo9Ckv1sfVkus/9lAFhMYxVLw6dVeHyDUiJSd4z7
HcaJ1+jRC6O+xUEPJ/T8hR5Fc7K7ggK05i/yNustYAiC84vpxG+fxM/3Bj+i4yjXXd+JoxcvsXeu
LeO3kRGDu9OFF2tKoc7OtNDbcxsgHCu5lwi2Z+vBYvr8kuCKTf3Qgy8VHczuHbFMcLEY9AIk0hJ2
sLmDWrMjWzFRIuXFO+ArrJ6Hh6oc5/AJ8HDymWH50FbTu7WeyEJM2yUsOgJl7ckdWBmolEEFSAFM
Ov6m7/tjkSninB8KWQUNOJeTFXlwkZ6HYsLqzkC3f8zGLCtOI4AzDp4mhmpc915eroZRurhAjBlF
kPGfLvd3oEyvFUIjzGAdhTKOpDuvMHgJoYRkx+hN800XfHLU5r/QuZjMir1jdo2QUqAVv/51u919
3kB8zcIjzMZgUA+rSj9h2H/DeoVIGnGw4bFfyolJ+DgfV/ekIIhm9Oi3HVYZir/FpZD6WzRU+kKe
0B+3Io/foXzOwYEI6LATm7LEYiLI+vOwAUNAcKYs/E5JIb/C4wi8bCeGCLMyHFBV6f7W8ci1Mnuz
tZo93Iya68ui+3cgJpyZWn3Z3P5nxE3DSZ3YSEJERudtHW44ekrVTDMZ1nIU67qWBUe2EuwPNUAF
rWBndKUcRcAv1dkNqpGw0dKaXWlQOujUnzplytjR59ISAuOcQKvRjEyAPR92lVD+4Pi0TpJyxQ9Y
i+QKjMhxCa7+0a8BpSt3cnuhw3WAArgEoJcBAmg0qxs0tR0d88J9++Qd/BtBOty25Hv5dTuvfI8l
O5wTpLmJmYXhxpDodgmj5wknq5wsNVhFHeV/S7zCycZrE3KAwkGHrH6U8nBUGMKZaWgpuvGSWHaB
smWHfqjaegBcKg568zjHkOfPkHnb37q2zg+A4ekxfR+AHtg+qWrjSbv91RYnMuDz0WJn15Bc/Fbo
VvbHheHvXygzS1QzLRIrE4leHF0/dRyRZ4BLefPVkFJBGxkbmj7U4htLLdL4wK9ycYNF3HoY1Tqy
bP8qVlM0eo/N/eEBp2GnHtdrldu4Vart33chPRCbhzeb7bWRw2UYrm0r5iyFiP/Et6QOwUcxkR4W
+lbzzPOMgpHzqMCO8Voab+oOMA0yh+Er/oKRZotE8bxYBVzzMJ00bCx6F4/dttgxv1IKHfc17f35
cE0xeIklc/PZFPN1homUtSu3fECebciS/ilTHFBhfTLOsP54F/CuncEsLQE4juoO0jsoOOG04kIy
9rzIhEKt48UY3WbAzlUOWis33eIzW47JKvoB+fLSyteIrCfHETApDMdekp6oJd5hCAbKhzK+lkK1
P61P+vi4B+xY5Az0ykfSeGx3za9FQkEyztdWkqRlnqWQjK/9WX8rV9VSfxDUquQPhR8gGdLKq2kI
MbQOqK0SqfTNfD0tQ+uSTsmBSO2cgckYK17s9Uf4rGMXf4xRVAhIlWn7xOtiWePU73h0Q/nQZMrX
Xs1503nmlS2dW7y6o3reuFNg1GlwfqlP8obaMarAw1enF2kzL/BO2aidtVHEesLztRf1UMrIjkC5
B8umSvLlCg2f/Jyzrw+fAMdtrmqrVlHY1iJbPu61T/XDnEOTwsxcTPcL/xu1aCMrRH98y6EeMxPq
goA4r9QCYUYNPTFfCxV9INesqQevUrXgw4VsyXHMCMdZFIQ/J66iN0K0KjekQDxi539nrAsUPCzP
8YZb79RTPbvH2gortFiOZjib8ZLA1BOC7+WbCnnfHWYSN5Mt+aP59wIRWtfSTMDVCoV4+kjKvhPQ
Hta5gNbzx1i5Wq8rirnRVVY6C47Sug452unZbjxEn3Kt7NEtPUNGWfURqQgObb0NFHT+/k4ShyjM
+ftsiKsI+zWbVwva/Z1wJt5ReBz6vYLLJab1uHDSTTN0G7WpFuoh3DowWK/tluUA2or1P4hpVbP7
zqAAVLOAYw4b0QBpvwTJE0pezfVQnBCT3iLnIU3yj8q3kh58hqFxu9WerivrwMGYZ99kq9H6ESRw
KaRrVSzJOxvHAKU3oGL2/zP/MLwR01ck0ES5lPM6jlQEweYGJATXbGOJuD1HfZ4w1LjRcAfsr7KQ
klZSZ3F2UhV2/lSb7iA0D5JVRg+OU7xlUWY1ICn+l0CJ86Fkjr6t4jIsVIigoTteAki1eDCGx7ou
2IXOVLK6bZx3Uw/va8Gb3ymyX/NEehXExxyo09sY0SdbLIjLk8vXo0Df6qLqRwa2dabxp+b72XZ8
/EG69rOTcJ3Xftu9pXrL2YdiQvwMqHx+rBL3H5kuVzMhFllSkJytqsF6Q/NiP8kJ5YVpm3oTvrRy
VKS5UdSMp+k4bv9EKFqIbXxPL8Wx3JkYsAmTtdpf3hA+UVOicFoVDYjiviKL5/Me/vk9BYoVLpS+
+TUCco0VrVDRW0QLAl+96Ay3Cme49YjtFe9JSzLVkHElx73TFIoFlw0gbw/OMQ6MgcXg/HFufIyP
lWSvXymszngNCsyqNqVoQReftLczveNqksGCAusEQ+8elNO3zMnENnqfzUwgivKworNIR1G4jTzZ
jww0mtAJGooA8LjD7qq9hXsWibrBvMLIQTt5jhWWxz4+d4dg5ph9l1bIeQ/nmWPSH3DBMgIgdKNm
k5a0/qqr0CHizK+biyYBp2z+l/pw3J7LRvgmbsOz7AamC8SPfgWih1iNnHc6e4FPc9r2p1Ktlr/0
6+rDr196qrdMnoS/i6vydw3r7chX3pZvzobn5gHWoEWIVaBg1maQQZEDGQ4R+H9OZ1VNW/+NwNal
oXnmwRiLagX9F9A6YTc5DuTFe/anLkzQ9wWZFTrFNX8zTM2lD7yXydZALriFH/PXmqpnBfhImhhf
T14sdqF5A43EkEv8b+fOcbbiM0q2130s4eUN3WhYBc0YyaYwAQEr/SBYgQlT8mWvLqgErjzNQaUp
MyiHcByXZiPHojNpIJ4qp52wcOxxN5lwTJKDulR6UAJ51cEbKzjGsnKhWPK3k+3cBdR7PvjOhyKx
ezKezL+4nvm7dzPicHnF3XO8fR+MBy34ZHxHLOHe3hH1AGUxGOm6T+NTHmlbFMozAbqBDMp1HfAA
+3aX8UJZpvKcOIhHtovNBThpIexauI3HaBj2i4vO+GMeFUrXXt2FY6jgB+uclwDiRV+z5L4nQBec
Ugd6XxyPrsCa874yRsHKOGi+WX+L3tJ01py10+BlAf0lg+lcXFttkE0DyG9FXhHnPWz5C91LDksP
lqdCfp+jy4DFZzLCaXCVciJfKOYddYwDOQgRnIqlHLcQfy91QSQa21TxWJ1iCzmbThmDD/gGqzBC
LOknBNapcDO1j3rxj15dI70aAuTMTEe8qSqnvXS7UU4f1u+dbVAGYum4YbPcoOo/S52L6v97ahdy
ykdF7phe2p16OphTP5FuFdOmQsu7IdLmKSZfPonqriAI9OsFZn9p5VG7vmjCtlgutWSRUoXALAQV
bMCYXNrwcDNhDFhiX+x5nDNtjw232GEpY4NbOGVlxQb+4c3sAsn0q6656PPRegxrNBdXSUeRfAK6
5scbUsreHtlskWIToPiTRBc7Yf6OINKNWL7hcd2t/jxVlBO+pO4r0bS+isl39uYzHGWK4U7l8K+S
0/WIbrEWerpH0r9ijQkDtyyfMtz2z5WhqoyYyyj4ML0rwY5ca9DQi5ad7FPKHvlZCtQEobjP6hQ+
Ua6IREfgTHTjLcqy7imEOD7OG5QrpvDTgRqfX3w3s1ujam5I5RzhoxmCntDksRyS6yVMQdtPkKyj
OpfHEHYFJp9r0XxAW3QMJDBcbVnFEeUmb1OiDj12GJw838m8f2whpMrdP89pGk8pESeLA/N7oRgE
lGhkQFBddJo7ZFFiA5a3O7Or5ecnYTPOgzKyIONjOnuQEIs5ELs4fPlKNM9W7dFEIzS4Vu0QGXFd
OxsZgSz41JAnyJ8/CPcpcfT2K6UhXALjwJJJEVzc5XJABpXrT11FmXgZlnkwy5d/lEYk13yypozU
nrV2ypx01cF7aueAXdRuOeDIGL5bPb6rl+4/FK0JJDpTDqapwE7Zcg88I8W30GqD0lFwGH1V8HVQ
xlspKplTY8WPJyPfxCEG1V0VoUosvCAoZDVqTxtIL1QwqqmTlucr73ejNdW+gyKSzPQTDYoUxsXR
OinwDFT1Vs70pQkMNYfeHD5MQdE+agI5i5Q6DnJ6qv6lSusOLkZq7zFOoryl0wg4JZs/t0s+IBRJ
7QfV4xKdHnQ9icHaPAk7mLYwhHahgzIzjpkRfZLQXpd8opV7G942Qs4tBDqY8KEB8+qZ2Y8NnaMW
Nod22GadIzd0Bo9cBKwOt+pzESO+iumFFVvB+517olVzp0s/1yPtQbQ/d9uofME+0T7ePm//zYQk
89RIBFDDiU6BcOO62hZ7JOHDLImDgg649G0iaLNQ9Z/JVj8KWL4bifTZcwGN7D+w+S+EcREIUBkV
LHH+9Zwpm7Gy2vU60/IbINHStyyS7JRy5UCaKk/Dg8YLYuzzsoBAml5juHfC66+6Hjylzd36gf1a
qPFTZ6UXgGblaBHA3uU4NQK/Lzc8kkz1nCN9G+fvG7KXl+Z5YEvSeDBuOrMxDlEpWB7WRYuOFlIR
sp4xWw6OgCVIhnGyzHkIHqwu8PDLpfLov7+X6OlvXhvGAaMAJzTExbFPvw3Ns3UPzThHwFkual3h
jl8tPXDGzDNYnl5XnQ4n1bD6+GLOIp5/YVRgtXPbvbvKr8NV00H7baPgJh+k2+dfXNC7A/SVDfC8
CyruQVqPi3+bK19JzxznQlkKdEAmX5F0dyCzrfNPlCqImm40ELITuv/3ft9GqL9e+WTWX9dA12jb
vczeu1fRCgBuYabB0aTAqllYk4FFZtMgPOkBNIfFyWhRBFJ0jOI7VDHqx35TbrLpNA16ZYRj8jPP
v7NSjQx6AImBfFzLKqAtDDEE3ffpu+6q1j3eOPVhsbFTgu2NkMBhzVIwykQ7uHs6UidllpJaxje0
cEyDQLEUbxf43tLIbLfpQfmrP2Qq7iK0RcJv9QDSeZVy94j+TxMxJx0zFB/Nfu6yvDhtedsDlHH6
79wSLubPaHANjjol46w4J5KV0hv2oJn2v7KfZiLPBgz/qjZtFGgJVGA1lz0JN3I+Lbtrua8q4+aC
fSbEyxdLkL8orHBAxJWXlLfFi1FfN4pyRHhc56xE8eV7gkiO08NUeg2gVAhAWe19MxKZdrYSG3Cd
vrTNw/t2E1/uaPYrNVF5Szx2+EMSxRSVG/Ntjn06XGuzN5Y155hHrvDNP0+uh6Bil49Q6nq0mnK9
kXzqGrdorQcpMBIkO6DKBixdyNkHOGT1E14Yks3RJTfRdjc4HC2ftAkkE/kMLc5XIPF4jidYzJDj
aHrdknP74926wUl+dy2u8h/kxgKVCb+n6tdBkVE2esyoVyLywYmv6K7yhYyeukjPlyxoTjjl6wDJ
j5wpNP8LAHUa/dElVuGjLn71Weao4AKeyCBB8rSlnzzV6Wbgoo09ZunzXPiu+VZtz4Ns91B/UeWB
2cS9ICRrz5BKcBT+Asn7f3YVV2Zv4U+2NNvTWrK8xWDjpcW9jLRdCgrlZ9KFRyJW6BWrITf2ZUME
PJpFZUwI8731tnucO/Wcuq3+2VNQZruLGQo3KxAnv4MHjTLj4+yAIhYOsy9plcXK8XjnNhb+ryig
QBU1zjHWjBhOlFxJt3LOZGxpV8Umulp6ZG8KhuHyN39sembp/Gov5+WPc/0Z/gu7iR+UvitXFjK0
jrom3BQ4dBdFxf8OanR3JD8NWjnVxauN7/BNLqw1BZsj/K4T2IhNL58Sfk7NWvWAqst/D1KnFRAn
kxswjvhWqn25/nzWpdY2xcdbaAyfIxnGx4CXUU0eMAWiwooKSDj0cels2G4shv7bje2XLfklk2q/
aVhdlxgudagR5/5UBzmlnUOoz/oVDpWLK9uLLIn/7V4wMcCK5uYNyfpIu/uDyAMyankAZLDUAK+P
EzqDAL1QQ82J2u8u7Ca7+/2FzA6aeuOqHY1ipV8AeqLILAyy1CuJC+Oxw/RyAkhHST5NfuMHw9OA
sF15eqtBbg3xjLDuHEuQFptepM7nIEFPEzil109wDg0g6Ep9KqsR9Kb48jMebeSv/i0ZzgBNk1aT
BK7wH/rKv0tgjII4bzQr4hXZfhNI+F4smgcO7L9YiNFVa6fr6+/EJsrIOxMgbLX55o3pDwJreHjz
Sfx2JPXQKNKs70y8QPLaFbr2LsCnE7RmHBG/VwayYUAJonGqbalpH3azeOqLBQPK7ALV3PW/jLGK
vsL8KE6/xjKlx49yCxuES5dWzOxCdj91EHuEQ0gXhR28XcMgYX/eFhM9qG3rnXrK4LHXuxpD1rjD
e3jkRCtQRRSJ29yhCQDMKYi3kVHyB6doCE351zsagefPzkbeKWvmgIhauMP0AUsuZxAOfQs0RPJ+
bNIqVvJ+GM3NV+lB/Da4n/0C5ZooTHDjIUBBJilVR6urG0Zhv5lZN0ifXus0ytW7bVc0KN2q0PVn
eeqyOnceZT9mTsnAy251KxOSX9dfXT7iSa7IrWK/0lAYacYGXyecY1uBYpyXWrSWwt0Jcf/EbdtC
zqQjJTVl5GEgND4jJ+aIWK5mijX5DJgQLIuXSO7zm5YHVCaPowVspchzqhFcr/Zu/CAsliUwbFhy
5vkj/FlcECJR2fscgpVegGNJv4bHnbTjM6PCTS4MgtXai6IJEScBIvTNR0e9slDJWcudoL6av2d0
pTASdNi763mNLE7rzi61xJMFxINzLd+F66eUjyfjWMlT27BYy8EjG1HvFnTmGc0whOzwozDrrJ5D
ROn7LDa2YoH5CnxLDb5ntvEQIYUGKS/aAMij2UubE+swPvNpts7U0GaE1EtTbEJBfOTr5vU1/KKu
J9V0/6VP4ab0nL5HnpIGABQkHuffGYViyv8NoaLhhDKx/OjSHNuN4U4RoT253BjNjN48w7lM/fhi
UjpnRjV6z+cocUN9YryYdPUfJXZGm8azZ9G9zbX7aQ0zU/Ma6KbU1grUdf1QyrgOpEHb/h+28gwg
r+ftt+B1XTHWOpib7pt8JXlfFtbZ+7jsuTmx2SW7Zrs+6fEEnafUbya4pWEghldWYXBAv6eoR0Ss
2fV38KoA+gb790DQsXPmFGrn3RvDdxpz0gs3ddJ/0W+ihyjKD+vdfsuU87Pz1WnZu6tAPdkXTLFt
oPor+IPMFLJsP5PgLdVLyJpfik0m5qFezxdCMW6QbDUTjAIESdZ+V+a1oR0MJPNfGExCYMeSNq12
mOpbI5FWgJ36VMyLQIn/0VsvpNVyKFJrUld+ePO2phnULOabdtRtgsTGMU+lbXHMB2XnKS4kO+Pe
DuJvQg31f+htIr445ojhFS8lv8idMkr4F4Wbax9/GgaZcDc1L7PGZ/GHonnFbRyKuMH9mMme2yuD
+ZczuHVz9/QqqGEG/4L+6/hPVdBlYH9crnTG0mIbZgKM//S/upVPzboTAbX3GfXIJxpwi9kxmqPP
/BgoxxCmby2wAK+jN9hBwfRaIaxnB78UWAtvdw9Wi5/fYXNFLZ7V0EMgsiqvnsMUykAsO8fU9sYR
kijqISGH2m7eoG5fApF/5LDc0aefX2mWIYsbkw78YE5XWQZhc5wjPigGxzbyJCeJ2+fL+/7Tb3NO
i3df5MK/0cPR6mjrHBRypD0681i22OoN4s/f1x2zloKjxBf1xL7jfCvGOpbJtvJEElMntZOB8i0I
9zxTfnqStPyh9gzKl3FmHAja9XHO6l5RIYnnfAgWi/wW8dBTqm0aCqfCXG0W9AIGeZSjT2nN7meX
n0ix3d7jWNJXgBL596DlNzVVARvRcujujp2PFpgWu599rDQVfgg7OY64SgnQ36XtWMpRY0v0JKi0
3D0jWBrEjvfd2Rg0MaILXRvgP9nE6N4ZCJhKGZ18qJP5HW/yH11+v+cJSoR0w83Wfv2UiJwaagjl
8/U6pDYteZb+DPJxq1Q2KW4v3NMTR0jr+fap4V5iMEA7B3zpKOeE3DEHqFIv6+Plyay87xNDHYro
eK4kN5cQw5821CSX1ea20wylLmeA8K6h5NMYlyIZnVGQCgECkNTsbLWpIHi/P1YyrzilICT9pZqf
oYqQKdboOYNMJ9QW9gd5P2V/EtEXVkZMhdvMf5nvfCzDbp7kIQTkDAYEfkpQz8JbyDeR/++geSix
GoTK6hK9ODRamMHc4afIGQNb/0RexhNu7VTt4IUV3YaDjSov4v2dpattn4bIyLfOGddyT4LbHcwN
bVj8UZJbGKTE+ZAaN9AHYPmt9s8eCcKPSsTVBW4q9lBXrPG2LVDIaTibL/9P8XJvngYBU/GhOX3S
Ts8ox5WZ2OPooL5KHydyv4a5HDjUGoap3aJdOQkmmDax8wyksjRIp+3xAe7Qh8P1+JEkotJfvxoy
+6kvkg9KMJGMh6cpqh+5H9mGQcbq69ufANymeapzKywhTHp2kGt7nncdT+Vb5yoRwgOtWpdrM0Lx
+tcSt/0ZCaR6opNX1VVVJ2R0KrZJKvu1z3B3e+Pm/eEVzM6VxxQS5anum+tYXGUKQ3YtzqSWIpPy
VLcKOtW+saI+b0p55Vlv5WlWuKj3Tf4ahFfTtgngssZ0MoywmdWU/77IgArSUOKIMa2O85VTSlwY
pvZ3SI7UHDtsXN3N4ligQfjS4cBbwjmFRhkwLi4tVmRPq9/9mI7iaJJjoJPHS7vY4dwMH/PHqvkH
gGgj6XqvclIuUb6uLmzo7Gg8qFOGJKuDJy6JiirGUUEiBL+St3FevibsC592kKh4hLkURi0pyHnB
uGy1cESo0Y9n+4DErV9mPuBe8YiF3W8LcEqfu+3DSi9DOeRAtFYDyu3gKDukqguE9Q07lMwpD9ij
WiTXhfK6LeznvG+eJhXlOJ4EtyRImX8eyauV8UwMNyQSvZTJ3X7d9kChbMQcV1DyVtAo7VDWflXz
cFsw5BcRWokgnLeYS4GwiGaKl699jk5lV3SKGj+ljz+ZE9s0ZRa/vPxfqzpu3Orcoz6Yt0JzzhnB
ose9Ccm2giOaHQ2Ix37Cucr5T2OJR/nPS2LIlQmhvOIdYp1WXMedG4T01I7/7BybMw5Oyu1gJ/Tr
MjRQe8d/NdtV7M1CF6gPY6GGCoeK6SXVEvJAH6L14Hyy9e6LKdIvWWTkk9ZZRGPqr6dAC3PdOy1p
+ofmIbd2U3+UQqo/Nv9uDgrxOS36i3y4Lq92UXhIsnetpNtmW3Bb+n2IAk1tAzGBQknZlnVf6iYQ
k8ix1XAlEKlGmjcdEM9USocahrb4dgXjgzUyp4y/5ixBQJaJ6TVMuN2gPsqseg2TpA6h1/m3ve4g
T1jyilNW9cSQ+WXOfLxDSPr2IQZ60XOVzqB3lSSzLlFcOk6wvhbeb6GjsSNZINQ/xnzkRqnYYopa
uaCv0E0ExzN3ExTwEOpj+PPjM7+DbA8gqNP3h6s4MV8rlbu+rjLGHpvJWkzjK4rFJTuXgzjlfuWx
UymKd+8/Ly8sTmbqxscg/LEvaZaBNLQCPOM9anbvRCSR0eQRn7F15oQF2D1yWUgnx6rXfplaNKN8
OirC/9TsL66lN9bkCLuyLPeiKrhUXKVwWtMpqlTwd6tcDoja2VKuIA+lAS35Cdr+Iw0zu/JIUJnB
+qQHeFmm/B7zBuxJcrEF0Y0QF0I+nHwcFxAT94/N+7FDuL/4FnNGIw+7Pfk8RHOqzcA+Gy5yfMOt
YFZ7Rq1ilcGqFniYzidSBAim7BjGLWEo0hVkCy68iSTuyh0DGRE9nuVKh4QUAOd2zqyDRnt3+Dn+
qMNgZe3uBuHyC/zfgVNYG4qO6dFQP4bl/dQ3Jc0GlQDcA2f/AvMeFEdxCvxU8wiQBHLwaRxTuiuv
ag9aYp5zS/1KbJ4QYYyQwJOaPB2d+KFM1RCOJ1rsAs4XMOKLboDYq/sQqaDCK91jMDRMqOtMnd+2
DVmSKQTAGS8WMubXDMf454fhLseSRYTwltjSOe+mJ80Zli5FuhEYd2fLSbRap94qWTU8R+FKhy4m
ToQ9AInZ2e4WAscsXYLxcJxI0yI4j2Hr2Om7pGtN7+KxFS9VB4uulXiguOz7lBF/+anYMCbPFul8
ph3DzbrRoXzQbNuZNi7ZpfluIK4aoXDi2KB7zY8ZzGHV2Ng7UpEGrZdg0HL3F6pqh5Tc0EWDCcqh
UbSFGQESMXu5NYf3kEISmHsCyUXMh8c/w0dATpr8P5NKb1sSIuWbhuVmBsnvtBOMOmXnXjG0DXNL
0pCnveSSuBMu9BcXvOiRg3DZzg5nDq8NJN3c3uSh5y+YTESvKvBB4gKF2Smlw1kzNSmUhyXqq4aa
YmrPUfepUjgqFt3CFEYwjny3nW/Lo9OcNfbvRToHj+g0h/m9Mkj4Ei0/lB5UTASgg5YcbNdM1b0B
ucGmrPEySYn9yDST9H0hHhcuowYYJteFFkYL1bsGAewMF+6/BHIcTXLtG184PpzXKrF0bWyRTaI3
7RPnfUvTTSuZTwwObptpc3Z+amJ9Eep4k14CXwcO6eBzJXgMtKBuNQxXQ+IxeA/0IGi7KfbkAj4s
8EpujiyL7fl5h8avt5SRbuqn8cHeRjnhbtNYT7awxXlqqQfDmsyNsj+aE0AUITp0TkAUjiucfvw+
Vlxitw/EkbYJ343iZwcAmOKIVP6FssNxvmuA3I4lkKtvzU8wsOiy5wvIMa3a7GPgRePhDefSGsrW
+WA5eJVoGwjXzQifSl5XabLcWAoURbgbaa8Wl/1unP8HNkKlR6kJp60tBHAC4zm4e2X6mdDR7M5a
K3MsMi97vFfgVuG+9nq0c5ME5WXDQJ4i/denKKGgTXbUPHmja9qJzcNRUGmN74Gd6EEAwTfrjS+r
qLyxi7/dKaIDSnGygF9LP8uFlhJVldbsOlwD9CwszXiOg10bNZeAnT5u42SWaxzC01KnxAUatRuR
xOz41NFdNytQQspbHrqBrmliEyxRKui6+6PNQ1eerWD9+OMwkpberwnA9gX8hqjEeFYVYBVA9PU8
eKbxNnkVjfcsyTObdZyDdnUfYf7FnE4ESWA4fQae+KX0eextk/ycfL1YIPM7r3Kopb1Gxzuk4f/j
RIRI8y+cnGKOHAIeDaHSN8OZPWMToJVS6wMAqoZXIgqWI2Hp8wiDqbqAj6PSUrOTBSHaX/Ghl1lm
CkN7cs4VPeU88QfN/xDsn0cOsD/ZAvm6LcNPqjIrkoAYOWYP4vlvx0OZadu7D4cV3mJZbP1fq03b
ACA0X8sNTQYhTF5lPtafiNBB8sqkBx8UnD6ZEAs+bKJMeKrZu8yl7AE+Q1lNqYa2IJ1ndLHIyEnr
vw0kh7Ocih1EWOGQRyacMyW2ektmdOzl/pPtVIpo6vym5h6e/ffqbwZG8eu0zGxVH5HGXdBTSRwS
5vIAT0JgNGS9GrEOBedUqRMkI9FZCbfTnQ41bOhTLSvuCyE7WhnTHSUGpK6ZxK5sO0bfT2JsrJpT
3+BhBiHm+vAOH579Rs4FlkIJCGFk88uUV6ebqJoK1rG2c6tLi9QZa7aoeOSqc24oWbaMC4LExsV6
JeAPyrxu8JlovirQ48MUHNqgKjenUM8ChqE/wIl1II3zoqLYIvsZ6yrFBqRnX3jpvX+wMflFRXGE
DfTtyusKK2kdZvnH4RZBvcUjKabGrVPa/qRuw/vbdzAus4d9m754qRo1R1C7JeFGXnz4nbvr+XtQ
6g6m6jFCZfiJmCTvCObTauKhtvQt2nRL10g28uWvjR9mcfp1b45s9SVrMAK8QqdoZbg5k41IHSjf
qrtli9UWNRaeITt+fXG1FAm/JBdQ1O166ivcQBcveTiCy2tM/coMWSQhAR+MOyGN4ZoXhFioc8yQ
ouspjTaXc77xeuKlxSVrDkboAnSxtP8R5a/lci1Bjam96Bac8d2y4wILJ5Ue6618Rv1qkYpzdsjx
uNnSwsuaz/iwORDm7zv8k5JacUxlICUUQ5Z4btcmn4sl/G2CVdDmHwRQszd2n5yb3ttdgaFl3M1r
nKyyAKPpR4Xr722beptJuesNtgOiL99gTvKp8J+gu7MYNoOFbWRbJO8JJ4zdXPOZJCN2VCm3GOH6
T3x4GTNeBrwXtIeCahNkSJ9hAoM5pipgF1Xmfm8vJ9kftO6ilngawfb55AJ4nCaLGxtRC48+l9m6
JPRR6nZKD/9ZwExCyhxO+HLuM/HPpWwxLrlbfBXpZLJrfEpC9OQ7sH927+mS0DNc5+rCijX8g3qJ
Ve1GWNNAv4ltg5Wjl4kHP+c/q1YMpLseDZpzVjTWbkWRnoI061FRRXWlBdafNAbsAnmFLlO+5ERI
g3uxn7a7f/j0mBQom59zmDGIAs1bTic8f/XTxKyfvnqc6yi98IircWLpUHdIkUbErXik2bR/vKSw
6YuYqw7JlA1Qgg3WMFgyPRDNieV60ZLCw2+kV1Ylw1UX/11HSZIuCh6J31Kt41ch+Z0tKmYOlmpB
mEIkkK5fs4Pw4JhBPkir+aBGoA9vmjgwAxv0ZjIcsMdg03k2S9oQGbLvEDV7OQqL70fVzNCwffvR
YixF3qalb+hCaW4GYjbesnFhuUkf75rch4HcBxS4s908bPzwZWkJ/VEWyKG1MbCjBvAJ4eVQMNnO
BhPBay4CE1TbJ/Yy6nDsQrcx9BTmpAvyGv87XOW190KYOR409wWjWYAxBd+NgGmKHApCXB/VMthL
hDB/KwPTiFBRyHX21b1avq7fu+8op2CDylAghAmH1L3DpVloZQMz+FxISZNpRflyQ/+fEIdjprXt
kmF9XOywBAlRLdnxrbYdmeLuPdrEimXVkcLZDUEfl4hvOf0djr04i2Zc1SZNRKo18eWn3z5xPLXG
38i0rjOn3BeppsomM+MB0eLv+LPX1wwGVYthd8BGpNFnmnyLGr5bf2gOS+BKSXODafewvHTHONZJ
lHrkMFV2cCxqvwYyur716iIySwSttWZbhtS5PSvXM0ZYiYgTfa1HmjGSXwhPOZUgLnDXIauLrkwK
vqg+f+pDCF++BZFTkHb9CB5Szus6L8KtOmppsmx+uSoQscg4HBsohroWGCsWy6GtAVXFPguZDpyd
kO07/iGPZ0YnCJUcN4Xr2Hjsvm9o3WZRFrU5tQDUu61aY9ItgHeDaMdcHu5lUdI5xzNvD+0bkLRb
7Hni1CHzCr5fPjOqJugOBmHU8ZuJNaKQWxawFAGR7D0Ep+lvCElbxlfRh/dAEqlZMTCWeedyYcS/
MZysESTK+FuGqwE8sTwTR5H/47DjEIzciR22fZx1cmNiI2Ox00rUGdA+vGb9wGjkqg15Tw45Z0PY
Tz2Tt714crNtUVGFfvdy0bJFLyJekXUwKd+5fp7xYRcLP4dBUzIDmBFBLF/ajmRfqmnXu5X80GWy
/o4be7uMnsmztsh8q55yB8PUl7gQOJbNDjEWluoqmWIMCWi2pyVAL+2UcXZENYqyRbPxO8DZcVQv
NhhAvdS+M0gWfeGku5V+Fk/AME90C4YvgR1lNIrNH0ddmh6mxKivnrkZuYKyQotRTrBd1ULY/pUV
DxQIeC1zu50o49Otju3wyanH3AH2oEJmOBSJlpHQf8bvFs/+jEUQ+U9vLWQ63ejRyT373+/2aNcv
5890yHJaCXtLLtoMLWiJ+q8dx0Iu0/67D77ayxRlToXgB2H5gqOfJy0hG8kK+YE7lykIMLvX0s4n
ISqWr4MYVTBQZ5t+ioad76xSk6FXXSvO9u0fomZcA5wSXw3toQwZmJaQEbjoGw6+r0DyuK+quFOH
Xd2n/qpmkV3t+TbBBTvQTGvfhWTwsG3GJ6xmb6kwBCIAv2/Zg7nDcM/kby+MZQ945aRVGkULgLJG
r9b9TFWbK1XfyFND/9MfzcjtdeoBkEBEG5a3Pa5HjRXs+QnoV0OSaN7/MmpxpBEPOxULF3t+niWd
Y6e8mJCdiaQm1j4EX2b8GcZw1FFccB/KVYEcuKEkfciInBUfYkwYahe/xGwidvStDcxNpmAQcP1g
nrtcAWCH3txsQonFfyiUYssSrkcY+4dNmtkw23Xk++/lQvxnYgdjNx5GqrVTtrWRALmdbaw83blN
R1vWbQNxQzGy+61nDg5evzv/WjYzRjkidofoRgkTolkjUOy4S6YkOftPKu2sqFvXOQqXR4LNviHh
5Oi9sBsRWjQL03fFK2xRLP2prURkI8ze/MhUfrzbgkCjwDEJZKQRbpV3P3KMHvwN5f9DsNob6E++
FGsqmAPzHhT8nRbiaPZOsDB+gY7CrGlDZpC9l/9zBFCe2ccD1bb0DSyDXDLPho94pIyijG7FXa3J
Bw8XHYyk9Xqp3gmUabRY/R2FXGeW64+u7UHicExZIRwi0bV5VJt1rnJ4+KQyn2R5x07C+CduP7Pm
cI0yGsNbjYqzn2HumrrcU4isddAVsOjdFUVKMPaNUZNqnq7KyDs9ZJE1iELW1d4BzzwTaXTFcHfn
QTLYvC8YSdWOAVDkKeTQ4DHPaS9hiOaVZ4r6iHwOZyZL7kGQRXxwHA2xWJ+Owa7q/L3juA2eh8I+
0TNZA9Udx3hLnIEZ5R8dM6vgj/AEzKqyfz49qeTIH+czWFpMz6Re8RaCaanoM+cyKRM/agq3JZZ6
qhfS6xG1IsbXJw5BjxaqjpQOPV40X8oWzKVZVBJTbzzPFkOMelD64PZIE+Ws6arCrvYUeqs57i63
XYZSokvkwKQSKHGZu+OW1iZGMwHbZlul7ulDiZYXaKSuoeYWU0JfKmTUNx74bJijxPqfRvOkFgFJ
Yo3INTk+jDATSyTTXQr48kEdhuwb3WG7skC/cfO27DKH7Q30prq3w2YM6/q+fIIxSP4G2NZx/QzY
WIyBV+qkTxYHx7pFWO3AHpRtSzOQ0GcBcpD4k6d+Hkke54nKlIS9tbJU2qDM26MtQY1ur9fHjhA3
RwmNLdnU4Muo3/6V6qM65C9ACCbKx/khiP0aB892k1BJsGJB1s3E8K3kewEr0zBJA3go5SQ9cAxM
rga1hTw6QdaUlUjF3uneDSpb2WwoV/Xrns4duUaPdgZEduoiFcAGTplgrjnaUFzz79DDK4Ji+D3s
Fk3y+TGMjTDig2hWKKSZPajIJqn71b1U/IE06TACNU/PJXwrfJrF+2czQVo0VMOsltgqJGF3H6a5
L0YgpJOd+ykC8fcyXoE9IJ40jJxC6oQZ1eDex6OZ4VjvvMDTERh0Z3DQPTKs6cBQ7FsT0SF8cEll
rYNga/8ULytWGbza5QS0UORCZSFtAfLNsD2NNy/oq+tyjqbhyny7W5DHGeQNm1Zk5dJGomoiK9dr
y0Y49AIDr8VIc+FdcQRgeSyeBs9a5/v/duax1tylv4dNtwlHHbCj0aU3MR6g72jPTs3e/XUQWegX
sMyyJFFlwQbThrCjINv+rGEbE0Jjx4fquk8od3NnY2XQTI6nQ+zSoYcqHwfh6V/VmvQjujZCaJeD
E10PV25uKM2G46DDDBtzdV4knx1SU7NkTTucnwHhndUHr1+UDyIPnBV3CHeKmiiu1HSUPHJdeaxD
GJMGNzJol4geG+1/6DYni9CpTV+MKn3cc8klZztJoDq4G4reeWiVVbQTyMd9VD9+BeS4iFaqZD/7
LYRAuJnv4Lt+TJW9gvBK8GfGik7fTtiX3V5r26QPLA1FXlwO8XxACv2+QtKXwu327N6cMo9D2Nwr
XtxFwThlkUF1oW/+wWNMmCgFQrU/VeyYihx/9bzAMeqTBWlCefpoRPCotsiGgoWfzGY6tq0I77KQ
UOnrhRvIdH1VF+cccT0UrLGO3XYbyk4pe7g2ovukfOunDRjNIZARJTb5+FvjhLWHpGpEKDzMz8zJ
+4wT0GlMzRq26lhTggYAo8Nw8R8Urzbpjf3vhzryObOTGS9YYE/xkzaA0T6WM/5yjiGYN+aOFR0E
nr1JJj5Zkot0WcdP+RPB/5LQMZDJ+iE6MUV/MD0F+T/Gp4kWHZowr7cHva4xrXnHPLQxnRM5vaqS
pTbRk18hfiABv+7u5xG5wmRkQMB7SFh6LygUkaoIMzgTdy0zmxt7ifDi7Q+c4h5m5JAWX/auOtFv
3XDN6Vexnoq+YrAwowwnV226cMj4SVGSZFUkuy+1qB3iaozNwOHJQ81+/uOkmgi1mEya6IRGulnv
Zkj3YMB+E1oFoNdZFtPAs2GIXpq/REO4/ECoEqOg0k2qTHBiiXjLgyjkHoijybt5maYDJknODiwh
1K1ZvkZ6g7Ci0N/Kv3oBWQcEc4pM3nVBNXQEtVM9S5lgzB84HovFNttUU1cyjxowPU73vDSTYgw1
IqcF1udhrg37gNCTdv+pU4SkD0MCuOJKLWynHSiGxOTTEgSgjEV49MCnmVPW2Qs2Jz/FxAVbK1Xm
AiziBIVJr5Teo6IHjCkvVMVarUChATcuD7NO4LZ8ioY/wELy62Se0n4bk6riDYjNqVAWvyCzdNdV
3rI4Da06487lb3W8011eoCfi5ucnccZJ6V58iBYkVdO1AMkgXJc/Ff52eWKU7bCmk796YIn2mtQi
jzPlSYG11stcJ3MOTddyzQ7H8yFrTsfKHLmKBrD4lDkhoJNpfg7tl28Nh+aJ0OWnbk132znlQAAC
AuYIpWCCHNdslL+Wct2nUXSeXlfYi4rWIigMrNz/RD5rpdsBDa4IdDyrTZd1LbFWXBrma4vr4JVr
9fPT5hE2fNOlEmuB7zXBgpvurpQ9dLHXwyhiW4MPcvPt0g6iiBNkGJSwzdRPED9iGnFhaYUmEqRd
NC6VXV5DQ+qusRxP5/caY1EpCg1D6oOno3oMLKeDumum3QkdQNS6KlraF9LhxSkPEat4+VJCJA5C
5FIhb2q4VWZnW5+Y3PxiVmvmKxwJRnbzjZY6wsmO33zBMSQLw2Fj6zuOo5L2K6aq9aW9V4tSlJDj
XCt/z/ndBJOvg/hA7H1dqDtuQmONWFD/V+Aak7vHbdrFdVGKropod1k822iLQt3X6vZVlbWUm6fE
8IcFt9PJddY7y1MorrwBldt7Vx8FiK/zWN8SNBHLADHtFy/fsXTn1USOfC0P/HfyGPYRVTd1mQCE
lMD6p4rahf3ijZWct5OQcfhQQqEcYY4RhSnq+U7HzeOI7kCkhJaXa/yXF9OJtVk/OYv/4XWcFA49
swT0IZeSfKKHXo8wjnfZXkXflriFTcf/33n3mLBwBeUZ5OyDDOSKWjFdMEKqNQLupEQcN7IC3KUK
i/VfRYase0mZYjShUzAZRYUAi27HCj9/LVZWZGVngt8m0gUhAPzzTZlhF80wCVl6YY3qS7crG5ox
aCBazu1lol00TTADTa/egGqZcoWSB/4g4iTZsKDLY4Zy0Bx5bSOD3eO30fzuQneXyNCEgj3TzOut
U+K1pSB7zUiD/6+MfnA/h3wpwj6Z4Y9zX3Q+lIB+oi496x0xOWGCRM9Y2gtCq3P64xx+zDC5PwwM
uGOTAgCIf5BqeXZhn08bwhrvtVr1YcGLZ1DCkZE/eq4r/2/pDY8W0W9gRrB9FmSFc/ceWtat9zCY
DO4LU33BLMrh9KlYpoTxgHUNHUmRvPqVJCZQfDQAaeIm0hTuaeuvGMdcFvqSB3pMAibaNaMlzXd+
iqUQTmXnUBkZHsARNhdaTdPFTAtJRywGZrb7XfN5zCILwfWyjUbDrH2zGGngiTn9oS+XiNTtJr4W
CdfFsUErLDi4PggZsUA2u5EmcEAz0JolVBeiKB97UjTgvf94SKJKmzOHOtB9PY6tTRkbJBL/MAzH
E6sd3UE26Atc341t7AwHyUh3sfY2iDoZ0pBo0NYaoFJHe4xjYxrKE30QuM7EG4MWN/S2IBKnkR//
NAppfkqu1VCm1MHCwqzHQXFD4e2EWUWmnZ4C+gDVdJy4+5wg63kLH478GdfRCS2tQE7ZSBxP4a6W
TR0Pz6415GtngQhpxPV9ntmEWLf6Ilk8r6DDbDIa6iWGzKdTbNACNLXie5jg43JcJgH4A38YNR0f
wCg+IiXKNUI2MoptUwwCESQ2JNQhnHlZjfxJ9tKSrOd5FJRduikYy8SRZd3lMVkARcIRMuUSMgYN
e37d9aLJVNsdo+m44ylNbWwSPfO1DXhosxLs/GDEaAHSS59euOWmKeTZAf/nZQAOhn5n8dAO3D+W
autx0iB7b+fqyqOPsq/EV1cKhGbbSzG5BI2qq1PUCCywTIAik/3wstvlIod0f7q3siPbLqGmdLdu
RfVwMKbsuCGXw4lOlafhlJPYpbFEvH+sZeU+TUYSkO4ZtXvDjHDRG7IlB4BDPvgphY9Wz+X129oS
KOJnhcRD/xb28K32h9UDIgMefi724XJSVFWmOL6Kwsa2jizdH6oP3MMXp8KUdzrpywBks0c8MErv
jLqA++5CkGK1eAv7txHibNp9wjRlP+z3K6yvH2/KONiXcEN7Kok5he4cj9BH9acsc/2Bi3+grN6O
Bvv2CluuLlJHIO0lTfDtUcPbaI4VdVwlBM+sE+wC/0OfPw7s+/+qFvQH8afuAjVum1GwYuoVkcNH
naok8rGrmJfq7fFRVoK2mQOHNr3i7zNa+Mmxh7ZuK+RMrVC6BClBWMJgPpicdNAZdpES3llqEBrK
rKeM9MHgyYXGCpV9oq1OtQMsC1o1IHw5mkCf+aJ4JBaqrRwKCLU0rHMsyIIiJ8MHjUMjHCtrZRTv
sqMua2ypsYQsk4OJZDuG2JZf3MA703loVZsjxGjP8QjZ+6OqVFnFzg0QjEgHd/SIxTgTm87ZWOLD
8Vo1i96+J7fo3crDEVviurRit9BQhuowS5fDvXYsx9hWbt41iZOc0qdSsMvsvHwN+vSIT0G33XUY
EjZXU1QJ23JBv0q4TgwThZwSS9TIo29IbS21WsJdP2td3DNKFbCaM/+CEHPJzdEK+yOW2pw4XMdZ
2DLQf/TsOkaOhVflqrnwmUegK8fKSecKyuqu1cZp5cGWDFvqik91J4a9c1ntylix12alTsjoFGXv
GmKLWmhLut324cwqCKH6on41WXWy8aBDOg80Fma2kIaOePH80E0YC3CUKTw0FGLsLo0WDF7A9MSK
8NuoP2coTW3EuQ83GZNlRJbw1e38NbhHXmd3XEet+ctMJfFOFCNb0JhBU9r7DafbB3MbRBp2hMCT
NwQgx6F1mSIBnqqtA4XGvHmIL10HoLDv6QOg+sypd0x8PhDvdUs8e2je+pb39tfop4FmGX/p9q91
ha+QneXIjyoJu6ioM+gTRAZN9eQR2cRtuXC5nGv4YrhyygOijhP6L/lrh6ORQhTs1QrG8UuWVH0M
dB1/N5F9r41yk2aA5ZgMzL5SAaSWVOV6qU4qnvblvLsz/q/cB1P3QxP/dFbjNIy1Qi9N/iN5cywb
1UndAaTMHzS25+O6LXHYpX+sCooP8gZ3SfTiDC1NhgBKfmkNX+osFN5XF3LIWRzsQZPsRSqEBEu2
NYaKgp7yM/NIQA+fYA8RIlArsUv2/5adXMfRnFgKw5Cque0Ng2YTjMZmSblgS9QxOiFNUSG592tx
bmDJycg+29qWrzdD2WmpmlG3Lzwer9wBh/XXZCUKUDvAGcamZfDTXpmzzKIul0jzNsGO60xZIdMt
ka40j5mEw3gZcQt704a6D5NiCdlI3eB1uQhZWXLJAyuPrhtbcKKi3U+qiCj3Tki/O2HfWBugbpZl
o4eXEst2j/SnbG0czEIlXUmphnVmcWwi5N5UyN96ahwwMc3mp82H5rFxDdka3KPZW81mVWqFglQN
A0lQkk5IePPQF3TTzPDJ0d22LS7BBJOuiQqCXHRf7+PTHIM9QF+BYEFvtuG0QjMwSyxv8vTyCAx7
ai0fAIHnyBss1WWkpwiIoEWBUGEOm9dQWS/yDUqQmbPBCgKzCpnTkh1CLhiCC0xHMMjr1AWrG12Y
HihEaZ04EBsf7ky0SX+cNUY0VYG5hiCKN0sNwRnZfb0JKDK6DWT/mGIlV1Uxc+wwgJ/5UQcn7qAy
S6jh8bWSYUtju2urbJgLUnojZfZSMqA5cmZHzCxgYaCau2WavQRAyqVh9KwblI6IXR9HK1stbdHZ
7BJXuGd57CI6mHgn98hpR5PLL1+u59t8XB0tCl/69cKEc/1Eha5beoXGQkST4nRdvx3woHcwxFmE
N3fP9uOLUmXrEf3jCyHMPxraPPa4uC9pQ1uDhrUJUf+ekEJ52RKA+gDLn/uwqKhQEgcvzspl1mFo
2inl4kPdjNoylTtP2havwIsuJWa4NOjVyBmiw3Ymb9LA6koRnaFYL7lv2FhXZxJDmi5A0U4nAVzg
MnHtcggwtjWahPzysSfcAXTktxaZ6aEjPSWVg5Zv0koQn8AiEGkw/zCzvafI9ObRUNNbos2yDMd/
EheB5LgoqPXErHP7wck59GIsdfEX1ZfMCkGO3na0NAsbnwKqczUVHg0RB8HRTLnvKGssdMdaCTqt
qjNK/Pog2wKVXimWz7JH0UJxSOrbBiJWSMVX2YcisweDXbzhC2vCfVkH4vG7hOZG8t8d6LZi7QRG
Stu1jKXzKtJIep0dPIDXsNSX0Z4SI8jB/KoOQgGysbCtBKKm3K6qgaYP4PdYJoK/bihM2H4EPvqO
W2+Z7KW/wyRkrmmRUPsqeVViou/5UgFrGW1QF+Ey90JuNqr/P+tQ+JgsaGemzQw25W1JxOp+IzMj
3M7xTkO1hsFcmqQtOoq1PI7FjPkBurPn05VmPfCgY3Nf1eMtsFukrsBNdZz66z5/QB/IhwuLz6Be
1cw90WTnBdHIsWefEPWFNyBxztQsTKku8UK5AQOCF7/JwudHz1eUPfXbbfeOlRRmMTv2e1xAAr9E
Sr/ctbpLDcip9iD4Rif7VrJ/7DwTKRO1CThEjHytM8My5iNAUvOoSMBa65P8sA08en3e2flekm6U
6wqfIXnB1cWcpUGeTlAzT5l/giUlLINhdzpICC1jNyMsgwzh+Txrt5xJUQceXdAWQXVJL2M0GDzb
vrGAb+vpDYeeoLSUlJLmSh4GgbCSdo+dgeYSXlrb3A8fgQ+gFG/OBfuIfowanBb7sBKOSAjuzhrl
PWy2YFNL9HsFYvKnzXweFfavEHT+wLrCUYzi6n7/Ve2MHuhPGFOTbwSw3J1CwhUZsyOCmZk17odj
9VcUwkgBFzIOcKXSZeMq3FAO04mgNiw+dU7muiV5/0u2f6zoPbsOqqqYlQGUO08cPnOXQrhKn30T
+NwFtYvfRcO2pstum6kJFUfEU2IBqScx5ytDgQd/vzd+lTbVtV6HBxrwgWjE+IN5+iVeqRN1OJKp
riSRr8h5DdzDVihH7of5ZIm2B+tth/YjuVW3TDXMBY2L1CmvBJhZI0dPuKRb7FhSZTyRQ0XfRRhc
iE3efhOMmFlFs/n16LBbSdzOm3MaGh8AeYrdIusrrCLPh8fOuLOn1ufzxZG7I45wL4Mdh/sdLMx7
cEVGyAbCQcf35Kgh5DoQ532V0qbfhQ0LJSa3JY8vmz09INtrfOI+I2XwgEmZz/XehFSYOvCOEqt9
tPgLcvN6iGJFbklxsmQHvYiScHfsxK0k6aTv0lPOk9QPSs4Fqzm3xFLQ/akJXBtweJXpUUUnR/wn
k5ybWinnHqx28tziKxdmLT9iijC7IpaziQ1azvUhXZVjNqdLqph9IrOHSFMO6inhJlG6GX+7Tl0C
9H36eDSnC9njfOJViy6bZlbgMjlGk5G8bPzQU3bkwM+BO4H01iq5wJqP5pfpARSmQh2cgDcIXyxu
ZWsvJMJaJCsuEgW8ytdTHdWB94K5C+wlNIW1WRcVs/FmUY623KwPHIB8bfv/Zjpn85qYKMqzn8QZ
+qnBZT0w+xjOReSLa72Fm39f7wdQdWxu4GL2ol1RJHKbrzTAEp7NRg4xRpQ+q9+2rIEE4MbZuMh9
XDfoCtCf+pTb5/PALba0JgQEn9q8Bzu1TiwKNmAiEa559T2vsSFgvjo0ujex9Y+N1Eidl/HR1cP4
dOv++Sn0HxvvfvsYo8cnFfd/rVAjZiC/b0BfRuYYOujYSb4nryaMM1urp7waCzEitdXBr5vhUT3k
XQOU3cRpVpTA2VMuDpveFuC/hAuuE6zjgZsr0TrXl6I9N1xz4TfHIpp7F5Z7OI6RX8xm2qhHfIJd
36/lnpjOys3jWEBufu32WgHEp8jk4ygQxbDT1DhJUkbOLr8Pqlz+PU+D3PmLkIM138c7mCKPtV9O
Aku55n2JwxTng0SZfOrjmViJ/vMSz/KnMXl9KtaHGk1KjqnUoWDDmo84uRn5rGcDtQ4vF7ACgbdD
XSxdXjePTbekC7YiGAdfApF00r28KUgpW9MRvo0EBk6p98l5qZl9o5M6obUm9y8SJwj7wavHw5t6
R7Lr4ZfF48uB2KEjT2+2RtCKEaUgVCAi4XG/fE6P/KEq0ibFhPzH0Y/BWt7D9q0uUdTzeuyhNd0o
K6/eYsN2hg7zsEPqkHNjydPYSMC5UJq7imTn4HLpiz1kvu1OHf1LOSGuig3Gs2NB88n8wBUvduOM
DkQn3mOPv26/gRzQUiGoxNNmroeGUQjyjCsvbUFCf1TMSNttD8sr8wix+QSwCDLZB3fox98n85gf
yyF0DQ4m1Z7C0ut9aXp47IpPCu2Xkpsf+ZYH6yeJ4vqaYz9W7WdBg/+rOF56RndbuxaEIlSI3fQ5
PfrJQTbYjX5JwDe2tL54UKOD1KmfVR6yYTPV/8nGDLYeu9p0MobQQtCqNS2bV9kwlfZj7zYlT/7a
MzJRsUpDI8PYA9aY+qru4M20mEVqxFKZ6hXAbFSE/6aOjyxBMAaXWlSx8pUGo4A6tTnGv8XnVzef
JUamBy52WLQMDgpMG9Arizqqc/mvWB7btYZYZimETfKzt0yWIc50yDeH0PwQkSwvyGrxuEU+xj6/
J2bFhKt42cxJdHU//ix4twO1xX6km0UzoMO1gtqwgDt+peOm41QZ9zzjsGE/FOxY6yrKPGlVLR0S
rQ/87Kxer5mAXMtAgRkMDbDtV4/1iGQHT+2ZsHuD+y0lsZof1VbhkvYHBBYRPg0qcEK4GbUgXoV8
xEQnhmpXQ53qSFZ9IMXSwXkDkJ3m7yvHo7Od/ctq3W2lDQNKuTR63ytYc8vU5hG7zyjYMo1DQBF9
uQJFynmxPrb8pvEz+09GYYPsic5op9/LQcYDPStnsjahUhmvQmxI+/z5swYHv/X+O0VZ0JBdE5k9
vrcFor5y1qTTtb8XcVebTa96IgIijZmVy/N4VO1Y9RnpTWuQ09Gl556Jve7dQwH1WGKEOotEmiXb
xWticFd+00Uyik/+saJ+82cQihUrAqYxq1Ri+hzCI/LbLNWeK1Sl/MdPpBTIH5Mn7o7YwgefBKkK
ditn33pL+h1HkiqV1H0h9sHwo4FuVwn9HpISjrMcF4MxCRnw67G3def7y71dzlKX1HSDrSVToN5V
ZyWPQFjntr5LKE92ZMXUOeiES/4waxFixUx1Fu2VkT/o/+7pTLxQ8ek1Kh0A/FFJ46wN6EjwOfed
pNDmdoNEFf7Cc4GUNdQOp1cY56OgzAafJY8/ukqPqSfnpNI0GywXd7qlHe0rjY+rMYnwjrFiBGz5
qNU8iUVLNnJlsnKjdUelYCZ2moXfWiCLZA/xGnU9lkymtGlx+KxqkS3IFWp2XMu3XeLq8+HKFIZE
PC7oNlk+Wp5x3IlsxpijZkPe3jaZQYP5xORt8hxJX4fm2TpsT/Ye2w1p/6lEI8STQuM9LkKKvxa8
ucF+f8f22cZFlan1ChDaz7qhkpI/1IBded0NxM8Vu7VVqoWTLa6QtfID+uzhh8E0jNx94oMFyXr0
gAyloJAvcgPv8ipYPgWGBNxVtJQF8GP6EZ5+Noxd5d1KCS+pN7ABBTMUDJwo0fGpjSmr9Iwrmq/E
LGQ7qBfquNRA6UDFoKE1nbezJpK1aBwRM7HMV79PAFYZ8Sel2zqF4tJd0Bc51CmWdtKwCCyJmk67
Zm3TtVuwPUgPWopFUguFOP5jcxQpfkdcWtq/0H/PSLTdmPYvQnaeuzTbBMuDV7z44FOj/MJuLORC
nkH7LM4GM2nYx+y98xxWTxvZFKw1FBn9hPBlHif9nOsrxOin7RD/T6GYkYBjw0vRKdGzhxCLhNFW
udxIQGUSNiWl4nVd3G2oHFV6FYioNM99RBRBwkTlQXopex8k91W47Pk9HuNsxW8XuCiLw+r0czmL
TXVIFGWrrFWpdluwj++ks+DN8Jmqpz+KTf+8QFf7rWmRfxR9WGtEF5+sGzJDEaJ0gqMQ4t1acVao
gXLuXojgFKvKeJ3SEROlO6zSfifm0ySLYFjKb+0q583o4UEEkbf4OiMGD3laakWoPpINMy/bgLik
n8ZqkJYmN09R56G4/WUwL5fawQM+H/+67R0e9SCQajHoZ+b7HZgigkfvlW8zRTEh7/ATujvzCUo1
mT+7gjiSTFQQzMYrqs2mo82hZP5XrHQfjHTQbpvq1eUj4itShXnvLMeAZ+x4oHUFJerBxioQHzh9
59ZPjXZcCl64T7eZYmNyrM0OnDoaCyLL+WDOSAeYfqLai5Gp72ohETUGXJRQjf1R1+Qke2a4uZLh
7RPpzHZqoQ3CwTx+5uTsYLJNzuc1dzgELwxY4jkPBBxQgh1//z0F+HMkcX7GLEVQxQ2FDvfr4yAn
aZk078qibnd3aaLNkwJHvyBfbYRjw81nmkdBaPaggOaNOqo8Ataf28MFWHVOvA1liNYwxANjIpi1
CssVFyTXjZJPpaB/abpXkTSe74hGqFazWOki0csl8w2ek0yt9HDXJvbJosKvc2LJo7TeRsAjkaAl
/XKJ26dvBwA2ACVzIng5GTc+Vm9L4pTQG47klczY7Q/KHHVbLcYqeSYURYKpfaI3WVuaaslQFGv0
QqcH0EV60NGKeIax9G9fC4SxiLbrg4MHxe4DXuL1P43gUXFlVWtNDtzuQzKQSo160ZITpd3OKdXU
vgs9N8knJP/HypGaGGGUjHtp15jXIJO0+YD/Ru5PMY6S8JRAFF2Gcrm9b/GP9d3fsXFJ2voVpaJX
vTaUwwqt7y2zLdWLVddhNScln0u/mBkDDlPzJAKBZCI2ag9Phs1D80Kul0muwdAikRVvd+YyB7jO
83vSQkFUl1+LM6qTYuG7C9Ds2GlltxgDmIEiv0C491fVtoVDfUTMArjwj3E9Wupt3E9oTjzX/+zk
pFx/6oa2gV9xUeXmNIbLxfRlSDS2kfqGvUwFVpRzYeu1E8uyWEyjY/6pmUmIUyrWjMhLYcEcHjwV
s75WThlAcS/c4yxHtJls93po1f1nlMUiCRlmYAw2octdR1bCn7g1b8sk/eZY7b3UOfeuS1Gf4oMu
otbNBSYdw8QpZAd1wPPesw7JvSQenYBF5m6q53Y11TZYl6f2qyZkI6OhWEbIMvnoC9FJFr5LRl+M
4KAyaP+aRgWTJrgJkEc75cOeee3zgs0Q6R2kZ/lQyRNSYoaIA+rqzIeUXh2QZk4SE1YkgXE6Ec0l
7WOCWsys0PpQZsnDcXNzNBCc3IQKVTYYm3WV1875BZUntBZUMHrYbUEJcplW2z2DKt7TdPHyD5jJ
UQK1hlsfICSrOZp/e1Ybl34sIAsM+jDCCxhTzbtxQXgPl33L2bczyJeyrCEWCWoeYwouVX/W3Nrq
HduMhGR741x1EwSDpWiT48NY9m8gRUDxOjtprrN1LsuXJfJymaxGca/2gfduG9d8+JaDWffP0JbS
xBL67KeEN18fMSiJJPwcqUYdZl7zc/G18deaXGs484Udyp41voOfjq+1D6VGwuuBXkRUQsmDn4Y4
jR+t9Ht9b+p/KINd2LpqnKqZwB54JkHIk+eFPaSeAs6Rhi6u5sABrfsGpHhnA0Y+speU+XRGrR2V
/+Z9sMIoaZW8dw/NMue//xDyfqAQitcJ1xgzu1e3tLuesbR+Dk5osRE2+y2ktqCX6VxKRQz7cJ7t
PFyxtJMcrT+E24NssVkuYFcP5fneobPqvyc4YpdXTzx8P/yGnvI/5IxxxdTM6hfBl6Pe0hFvS7qI
Nft744rTkBZywtjiml1M/CAUTc4018+IldU4F2ZL3SHziF449rF3RTswV60Yql7Hs+aHHAF6hqLS
KZOuXhKVeA+FadFgWKe6mxHrYvgwI08TfoHtzYqw3swOtcMXJ6Ip3/kftvzzsEe2vdWAFUfIBC6O
Gb9EHxakKGdXzDDv5jJq26PXDa0c/llPdXrexK3cA5+VELzduOH+9nYh3ytSl0lVF4MDPH8DKl/s
Jii4x2R15O6ouUEfINSt0tDI+aNwyUPPW+MTvWz7LOspR+RG9Uzp91zH0/kAkrJiosOoyWaphJDX
GSBjD9RwHLqRz8v9rvoo25S7oMWN4gfWyDfxTUEFh/4XxRMYxGYOC6glcW/rP5bLNrYX2MPNBeU4
eaJZAoRlq/tFZAGx60QfpdMOnr/kUAYY8ExoDt9maM2edGGz6vC2JfGhpHfsH5wZhslucqYL//Rp
YWEUDLkGTIfjAnD/sXxP9h4biqOooNJB5/5ewUyJ8ZWsRXX1FTkxQs4uX7URWNq5VA5/Wb8FbA2T
9b3s3+EPrR/clGeMXo2P8ckpy50gWq1NM0Qc0XX0l/Z78L3R0C19rQKTNmrVMhiBWYFqE3+e3PcD
MQZuQAlFuHBritqk++dXF83cjT3u1MQzSkgalXHeeXQk+buQflslc84QrMUv1hwR+F1AmsA7EAjg
Wn+tBnO4VYCvLqL6xxbkozLBnRdLQo8kSTsZcZZxSlP5rSgcVtNuWk6MG0hPRTPZFFralSjnX2N9
Zna6tLbwSDLiXgZTmYz++WxOJqO/5PHCyd+0bhWMOYZWZ6EeIlqBe+T+ljnB2U9BxArqiAcbum02
Zg3ngwG3KqD4Zgth1L2oC6E4CqJzmpBYeHQNR5XTr2bW8oqh+VS1nDzHo3X+09pixBzB8P0kaZLz
lpbcMdsgInsFpD3N6VHEqp0cHZ88Y0o+fZIQBu2N1iUorLM/A7ZpjCOesTo9z9j6968PurE1lkYE
FA+0vG0oWBVM71lnUXXs/auV7ZnBKai+Vk5Sg/SdeaCu0mjb3sfwkTsU257WXKeGJPbOnM5B2uvv
5g1nTZqITvLlzfCHkpf1Fi8IhJVknZO0p95z67x8tRtQYOk7gllBWmyvhL6ndJlik2VB1ayeZm1z
dd4bdlXFC1lESh0OCg1dlYKLhOGoUqhY+bA1gB4OxOM3Uj1jgEAXbDx1Wy2SvY+uWQNEUkR5lcYn
GKaGoMrFiulLTFVQ+Vdmdb3Bap8g5RbI9OnAxOqUIaBvOlcA4iOCHeEIguXzgI/suMFRqIShlvRk
GOpYEbHd+8cGm2PNm21IBaoife9RW6Nsqns2MBVnH0TxkQJVTgRzp5zp9LBuAgzKOhuk9smtOCqp
R+fZ2VvD66PKe6NcDzZIMpV8DbeDvdZTp+rD5rOKzeWUZUnLvJwoPYNjEiiPlumgfJxNO9+M2iDF
ofiCq4fT3nJbDX+w88Bj0K1rto8/+xmTDXX4mf8TGzVYMhmuDt1PSco1p/Oasso6PwKnvLkAy/92
yYkZuuN4eBXie3rUcDtN0ChmUq5gko1w5iM1R3T53qVLRsBNs2bv+vMBWvxq8C1kWhAXMQ1cBJdc
F9Q2u68V//4GJqr730+1t6xXPtKAdy1UyQVb1AS+vkK+NplwDJMjFdENgY4Fv3aLIWyu++cVzS2y
ODIJhppvKq+f6bzTo6s2f7D1JJnh0T6qy8r15MIzMC2XCv115eR+v+be/uUyj3s5qB6V54qIjjXp
JPrw++YDK875QIQ2KingYOw5hTupLyCApaVxkc6LuwOdMQlep6REncl4x/31krGbHVZKpCmr5L7F
X04D6RYIsE/l0bytpicw6c5qaKKG+Bm1ltKxTMxTHDX9oeXS1ygpf2k+qOSJ2PBRf2zsSAgLhskm
njHEGn94xjZCd35cJasRVdy+i9RemdVUr7/JIp81l2vuGTxrl/AoTf4/fAkBdXNQ6jX2oHiBzTFe
zfHDqPrLwax3I8dg/1r4MbV/aS8aFsPOFZK+KmrQWVDKikrpLlwDJ0gkIOWolOA4xHs7bDlfstrD
5eEOOx2Zf8fu3+H5+lOF+6OpgoVHpSTwixqPEGTZWak4V9me0X2a2BuRniDxkPmmkg9/WT3SFQyX
YuhGZGRqqxrbOkXM5067Cm6n5UEz8kh+dDzelIvezsIQViX3lXaSwJYQAUmGLehL/XR2NGrp7tDZ
/+6feA4FEioXCtRqXqT2MIP3K9IKl868qJBzZmRnZsLfwTgjTNtInHJPMI7j5xJW96kGT2WYUVKl
gtYSQwxJcVoQ67CS6iXs5JxvCddltXLidDOeVHJgGZsQUSnCA7hkFvjlDQ+fbXP7JaJlNUfKgLHB
vF7BgaFWjTkCWViQGshHNG9xFUNJ9kLfkf71v0t2P98fwpJMtjiMFFfTIjHpQLQjtTfkW6+vWaQ0
BW1UJ20y18D0xjDYdytRqcK5r+B0K0G+Lo+TDNulHx9Is50JL1X9Xfjzl7NpMbd5eRLjmVB5M56k
G0TypUEXGFpZMLhM79jkFsOmmuwb8OpdZzaO1qCcOBLFb/Y64snaB4EhP5ayA0Ynxyxbe6CqDzyQ
eiVVMZQZaZMBsm8wfocZ1qv/x1FH+nCVuQhmFpAwb70Q9vBVdgsJPoY0Q936UZgUun2hpAFtx4kk
cSvKrGRCPkbIaon2EOIlQFKf9cmg7S4ZG9RCq1C92/sk9yCUzLQ2ors/w9aWytdiDrEJWteiPgqn
YzfsEH6jxzFPTfBq73DFCfRVYUw/HiQoPeMKSX1KI1TJ8kziEVZU+9Sc4IDq1bO0KDpqxPFM1G++
62dbDKNA+PWuCTUpMUShlnv4aVMXgmb6kaJX8l/Dfx9mmap7nUg5G2C9U14g0OQjh6FX/6Czekaa
I/6d9/hW82wKVPjcDbujnDRZ6IjY9ASvD6q2ZDwku1nqYVvKYBaucX1itSAkhtItjocseJthcjqC
fLJdK9S3xm3iQVpWfi/wEr9rkBezFincHGPDx3rqUtWaTREbxQ0IMTrDNpiKQbkmMQAV3pqkRwnE
6dEEGySjDGPyQiBQA2+jrpQxSM6ZTdQ7ad+1BCh+Q9MCcUHbX6BCmKS0RofnwBnPCrsq8/bEoOpu
t8ojORL90v/Nova5pfUlotGJgWVVeOB5dKN+IjdN2uoySMPAc9BN40j5sQkq0cZnvdY/3b9KHGpK
MePqrpAc+e6c7s6lAF/ulharL58M/WU0pl7uO/gVrYRSfYZ2EXe6VEyuu/q+N2jrDFz6IHIWHENf
tDkkQKZwV9Ypw2HoJ50cCU8aubqCoI63YAbLT13zhG/MWPF/saktYOyTJ0U10nWIyPStY0xA8CIQ
er+C+IChpUgH4QlRPrfMjOFFcQEgLTbhDsyu0e67gZSWpsrqOkFloWXgOjuRGB8VuFpppww0hyL5
0uDSU3GIyu9y2EH26b/LSLCg6fF4F8f0EBQtX75hk2BUmv0GDht+67B0j+ekRtuPXp4zTCohHMPH
hy9IdVpNN0C3mTVOYm1Rn+7Bz7m1Mh4WD40xVEGAvoMiyyTwZel5/Z0lsf9Zdnn6XH7WlUnrdmsL
fTbVNM5FAZZwOU7oRKj25vbaO6QOVzjt8iJa5oBqceQBM3z9BZ3SxIvykV40G3+4lJyNbOKuGhdF
SdMeIGKFuFiPKofeLdovhdbpI0tCMrLfcjk/dfM1UligCFjeze3c4dGL1odUNsEzy57CdzkE/sS2
5OvbiVaEjimuVlW8/h+CdEVELbavUps1ULLMQPd25H1hNcr7Brz4teZ3InWUUfxfRDp4zIYrHoxw
IEao8AhaeC+GPF6HmBLAxuUkSf0z+XPcoCfd1Ab9jwRbCnbdc29VBMLrwVmUs6VMJCFuuN7Nmmev
3cpWk4oeb1XDFuFrdmhpmpDSWgnD//EIeFqi90wX8KtpM+T7KwFA0CA26dd2XH0yZ8tDWIdSBeRb
qy2FwiyXOLt2Mre0DaKOhtEQF2U54VSe6dpA9EwzgLEirMSqhsqepyZe4uqblFQg5it2PwcdWf/X
QxlDni7vIsMQSoHrtA8hxqSWqxXon6FnRlaisWM2JjqPwpaqo87ItMh4ZZgBJZHaoGgTejrfi+u8
b8biGNePpp505zBQTQfu/wEOyYRHY5jVY1Jv7k6MaPXPdEDoGx2JxInYtFE0zGmIxtYxNEc1AI8E
iCtw4X8zxFLczwKcpbV5NMWzeBH852pQDvfeKbGLDGurVQ2wtoY7ZuXh3jKgCJvjJrGpG8kYp3HB
l3QcfwIFO4R1IGSrWz5T/cJA7ADrVrjrtE+pDqyUU5ExOJVBAZl0k+V6GxrjTlfPRIKGzlmH9LrL
oI3IxwOzHks7ukl76IBZNSulXmrvX6gtwU/ewyTm0AL2QANvtl0zfVQH4GXYCvpRtoXFGbazIkJc
1B9NyFQYqa7Od+ytfVw0IHm44r3CLbRJdhPd9K6DD4DRLWhDa+nwt7VUFlFKybMe4eQhsLxob2Pm
G/0Tm9CituMNnOtIip6enArWmoswg3RGSXQWibNVUfIT/RFq9U5xdgY4tu+GxJ1I4R7xCSEGbQIm
j9ef+pq1bk7LlQGbkg4G9m+EUQE8hlcqvfGJQraNrkdeMAvbSYuuFj75XxtuRvU5FEu3Ts7TwUeG
9aGWh3VSS6NdnjhaCH9xr02bGp4kyeswIzSJ/bWRYWuWwrq70zy8S/ByTWgdYzbSyhTaOTwaf9D0
ISKnzt7/eE+nMgW/WYQlVnwe3cQViFqPxd/8RYXWNGcQsdjZmkBiY7InyYDol1ScfY7wlG4AIn88
+MRYR2yEwjC9jdk6KcgCD+vnwStx7qrAnLgYZ0AX8A0M0W9k8OSf1xgDntZ6kEgoB3aSfq5ykphK
D+9Vgr8CUpz/Y/YCDerx0I9NF7jRe1jXmBeTGfvzuGXkPow7ff8xSk2m6veFyRl9JEVpEBwygYfM
RcPGqHbBSkom8pY6ugNB8ZGAARpIlj8A0VKFPzFJePNOJcfckkh2Q1aGrzyzRaNudVAyNFSKGCIn
LlVUv8VdHQmLIswKRk3UA0/RYZMNSpisjwZ7lzsw1+K+Dj6mPzo1MtlmOyQf41ii2NWUpTqmREWt
to5xq31Gor7nWbJtAf9a6MkGnyL2N/rZJOk9khD0XjjCnpSX6122Xdd1CTNfyxiugXufElwAivEn
bFBXU1UcOYHUnmd6sXYIvVpfYLI6Cl9wdyFpz51j/KFPK6upvIj2Iue1gcSVOSrbjLty69Csv2/l
lDUHob5rNkkWb9Ox5maWjnS0QHKnXDF1vm2ClaeJ5T4rG6Tslbgmk/vwOqKa0bbU1WK29vKWzqQ5
65BUJVgfSiMO5wgHvAeXZe6HBpPiXKPES1UL0aSbyjx9mTyGoysuL05bMmQHlejg3oISY1Ls0Q5j
jNVo/o7teFRS6A7sxOruiC9fLXYYOnkjoZEQoGx1v0eW0bYrtF85vAY75hco5s0V5jyL7qiBATHS
c9B1PZ0Hd3iPDR2QPRbzzUblq8gPLUkwkrr+JWBrjmn8CPAzXFZ/DCOOjDGXfaMRNhLH0zehrpWj
75li/m4p1SSSpQfrEaAfgGaq7zjj3n/J0CzWuUmVYExJ22llsvWQ4LX6tEHOQnEVskO3IMFSkAdO
6q1PeM5yjSOOjyKA8yoGRG6YWAJNWi7jRlHIX19ybjVHWR5/uuYBaNfFzroLDJjdyF8ChiLEdTTt
uEyjLw5uNh6xYxLdQR1w162BMiwnQqbwyiwyZCYBeexEthlrqe9uejwznuzz8c5kJxtpoXExk5lS
Z71YdHNzaydfSmszB6nxxWSIBftU6cVeE6YPmdio/NQZMXFcs3LBjq5MOl94lUoci5NwQf5TXYjM
qVv12loHZtiBC3Eb2nnqZL1BpC6MHRqm2s0otykSA0MWkgDZ3ydhysIrO2FpBNyoxGz2usTgo957
65ddjVW1uK5iL5YgQsh97iXe+ZoCI5tPaFsXzeUoEFIQnwf2WC2+LCGR/inMMiTpGMuHFZB1j+4t
wJEAmYH6oAq8On01Bnnf5br4iFAl76pU6Ow8mlCvZGZUPNw1JqSb38eKtRJchum+xztU5poEvylx
gK+unRl2peq3ML96I96DV4Flk9sNDt64HwTObHb2S2shOnWj+LZy5u3p0KTtzNNBWQ6dkyRF/Ec2
tLWgw3qXhPKVovCL9YQRW/yeu9NRrbFWIyO6W41UbtQiGwksufzdk2tr97fM0aarygrj+xVL9Ot4
l7KjJaT3fIYbSFeNaZk0SNFH6QdkH4aUMdLwU/GAd/FU0ZuZd4si6Fz2pgs8dCEiwV9m8Aom4/8J
pO6lgqd6IoyVG2eKIucxLcWIivawdlz3Q2goxFkhvv7+sNrJudjVmlMdl07K9DxlrKSSYKOrFvJn
kfTB+BH12oYW7r2LRW3afGQkvWe4UCVbAYoc3062y/UNluVN+Dad8EpbhKgL+iqshTv1SpDvksSQ
cG+SguIDszvYIYwD0RTnUiBEoOGxnQGaotUprRpc4T2J9Muc1X7v87P/Dd2V0/Gt8pWcze4BJKUr
wOyndw3tHQKRy5zqBr7yxd1GBMQf/g74+7UqatupNfTxYWbOdW8QsQCJNoh4lvm5AmDUxaSvUWxJ
/nFO1upH5x+Zgpp2lQazgyKayXjXYkqHrawU23GWkEqPleUDUiCkzpsZJ8VBnHvITVVv1JJyaPa1
Eq8Qgs/wnFaxsrPAz7dAMxvz+E9fCSD6dCMdvFzg2cYq6SXLpxaP+2DkTADrIRht8Utn0e5pvrGC
bQb0GzTUDzHLn1ZctMMG1IE6rxY7zRJmGvazIqs0eqUtXLl0MPjBLMmS8VjBTtO5xD5VtX34W0sA
MKICsnsGDtOmrItEyAHxCL5S8fsh9G/MsoSNeoR4ejaWiQ1Pl136ZGNGBdHcMNnOfYHo0BNP4STU
0Tnu4bkVSF8txMnoA8zUkAsOiPsi3rB1XE9VPQ4D8SvJa1T4FJTU1TtN+bGv0YkWG+NtiGUFD1Kw
zB/rvJHuvhQNKzYthxAvVAJDpjEoFG2WwJz0A5514+eMF9AWRKeSSgFuj3QB10Z+LxyR5YvSHEia
lGaIbyXD2Rp2nROUIyE6IZdZ591OcQZHPB2IBrETGOp9SHJhbaVXeaHz3JI+yofTMrHbo+XR3w1g
fuZ7+qcJyKggk8OG3kCx21baX82UnDSsVJes6ZSCIsw/mt/lxxE/TxpVK1/7BcfdctWX3YjGzTYl
8hW8i9BQkRla3f9s50URnZ/vi3b3hkzm+OzthuaWlD8NM8kZCyCdIk6kLNESGarTZubplEPiLp4c
JDWD7bu5jC+mE4H4AhKgBoz5c6HHSfpcGYKLbThPcPIj6qXjiTALwJKCiSXLmb3tHBymXidk10VR
tVrrzkSpsjVMdqJClfggWiWsyZvMgb9PMxjRcPywbQ5M7W7ZZYamjW0dm2xTuZR3tL+1se3tadCw
JMtY5GyQE11msfFJozl/2p7IAWS+O0EgNxFuxa2+hRSMCBqg4khGMsHGlJOKFNWKB8icp84l2OVr
ZI3AOOn/LaR2WbJBvjYlWp/mKLOhsEiX5n3t3LcehSks41osOMGNcuQ3us2wLsLe8LvEpWuwXI5q
srm94IZcj4bNwL5AqQ0LgProOhajR47VMityaC2jkDcQEbrD5soBh2Ztah1FoV7tRQMOOpTfIohp
ZFFMeZ6Z3A26QOH0bKE02Kwu2FijkngdCqPNaKgPjHD3R7/jniGQOGGPzcSHNtmejQpJS7tV1xDr
5HBSdhMnClcPh3kLgFRK/WJfFwz6D/Q28PXz0juPdzcVbN4AGeejyz7CtJueNxXPmtcikhBBPVb5
NnyH/11+pzjWi3xHAT1y1+6yY3XOp6S7rbeytZ4CDt/0sUAAJ9nXpQHl5VK5WEgGk0BAoRLkxh2u
bYDZJTfotv9no4/F500EzyLMm8yMfql1v2+Zu3U5enztrdbQRjMYJwrwKC27rpboylBqwmlkchg9
irC694+vhQnQoqHw4fbAVU2WiqYzGoIaQYWGvU+6i1u+3xgsLOCZConvO8J9oWNDJfV/d1wg87/u
3UzLHBM4tfJrU6laUJZntjbOgGyPAcENHOcSSlIkVMg/jN6/iHVnKRfipXDnkx73Ef7MpfOmuuNG
PbngKzeAiwmKGOGKW7iGaCt+qTBLuEiV1QLIy/ca8Ra4zCoy9tE0e3bvJRpELf1wlP1t+nc6Fs7C
6i2cewlLkFDGYs4lNIpN2GNE8xa49REUO3lE+GOjk8gBMLlJz7pvo73dx1tX6six8/+SVQWbKso1
VpnHZRnunj7Act3/F2rJm5d8bRPh8UJG8nvADsFyILS4hXmbdnysChVFBDEaOgOGyFBabNSEA/ju
0EtLArcnMK1TrWW3KeK3rvSSWtoAZrPxAtmXWq7aA5tMyxogqzmB1BwE+6xBU+td1yBkJ+P3SgSQ
PVqXbEz437dOfNahMSRG+Ai54y5qqHO6rpJ+ELPJejMouWVhCIVW6Yd1VzuV+lZG26p3GmMiFiAg
YLtt/yfJunGLXmf/t1rSc2uC1slOPlO445W/Y4RjcPCGqJDtV8fEt+VzWsR8UZwR35mYFP5eF9lt
ekClzpLSjuEmriqHH8+gealYtIwPFA1tsfKjMZsHpF/7q0dvTe1oJ9BjfLlPmn0fBIWI9kLvGENP
cP6FOfmWy2MsZnBxrr2dxbTViY399G1IuG9KNvvY+9ztGbBi5KvIxpBG/ajlJzVsWhzsbpHARj07
l3KCwvS2VXb6/KokQIiRYTHHFaxnCNQ7lFC/WtXBCVVZgw1GspDjM0IHHGVNM0zdyDTid9e8Auzi
qLpTYAyqsvJKI4DAwqfcGurHNHy0M5RqTycXgaqITJ78S0LTjOHG+Aj/96yM/cUmuXiY9bzreYWf
4380wkYstMrJxh8SJCbynaj0+lNcT5jZm0cDJ43Up01Myh6b+z2ElSW0WOmjL7aIsZ1Gh/Jm48AS
01CFcDuxm9lbHrKZ/aPcs8mhmO3IBTA3oFh8wdZPFv56DeF6W1R4iw3AsGxIzAkLAAQnFkZGslxB
9XXiLF25gv2100nTBQW/611iQ2znWMpumEpWPFXQoZBNQJfLY+0YGpj8MWvAViAlltsXW/4cCZCJ
sjpjVtIcu/gIRlE8M2H3sHQdxvt9N6E34xbXTIdbI5yFJSIt5UVOPjbRHrwQukZCqzsyOcje7rIN
0SyTrmPEMaTckypWhQ/awq6Tl/hnaHXSm49gI7I87/Oc5l4BwJLhln6Muq2sXsuM3oDc2CPVKhuN
ij2JfjDs6197IFyOa7IDuRz7opJKUj0rKsbH5ygXSUFN4XFDO7bIpmXkiRUmtZuoEobsbUQ55n1X
6I3B5lQZ9auhkPUjz09LMTi/2xyl86Tu5X+L7IqvtML82LWppJbBko5PP5Et1T87WhBbiN5mMxQD
r3HWAlw+saW8dpib9ndToKsGMpKYRN8W1iK9+bCB78W0AEmAQRZFta4AqsLL90Yww759hpQerIeW
dq2JCA835vMYYj5eJweXelJRTwH20iUOqO395BdI/N/IdHRbHIJT72UPNsLfhzRrEKXx008G7420
Iuo5ApO6gJzccNGrpdvdDw1F2LvLF1UZATijrrsmkHBva6UmuZMB4OgjMxtyLOIbzo0aafAfYNsR
KOOfNOuFuDpz7A5O2hquUPNtoIHKEo9etVBvYP+uukxFKbjQ1Uojw/fxAHNOOKdLLhqXPReQLQ0B
Tr8Jb7Vm2SH/ZjGyR0+H6Kho9cpJrmVAMOkB2Vr/XMfxzvmoH4ynZb85+ChM26mfc3Jp6rZRqn0x
/+aH6eDdv9i/jmP1/X1+ZA2gjuGYXLury29mYJKmSyJrwxoD4rYaQNvmvNUpNt4FWRmcrPwqHL/Z
Vn72nDkpAaZNVWMs6uF4MQ+nOSS3Mc3gav0qCP+Z3WYONNKxzB2qn24dT3Z4HlPuSBQhEO6kBMFp
/O5UJ2x95CKLoeib7dbASj+6kXNzPS2KbNZF9vHaMdKc1YnkK0xNbBxEEt3U40UgT8CKni3LqrYj
tM/DjSAlL+R1QreTNhX5zZ/CXQOHUg+31Sa7CR6GCrSJB79pYVKEsZqULfrOV/rHZ5nT4JuWEzxd
O19qpJYo+0OgHak7BTPD8+SL//QiSad8qk328C3hKgqjSd0DjiVi/2iccLFrk6wsziAVIDB1KVvh
WiKPOJAYh3FgfVN8lTknMPMkDLghLiGNaQWXnE4/52Sr8HhWlbfFWHg8BDQDpxUtMOjfR7HK72pE
Z32RNiLQ9/PfbPVA3HAnGvSm4q+6qKYbgV8CB2wEK7Ygjk+PtwIgAshbtNgEGaU8dsXzvwbuuqit
d6Oce3DV4xJ1CLgdcmyqSC8ZGjTSM1bnmnhW6nFRE6r2ZKrPQGRJzrBNxm7PWickyngS3yYx/maB
WqPXB2NARCuts8qkTcNWikoLi07yIYhnGB/My7UrBAaZnef9K5vxSd+P/GkqVUQKf3wjXA6GvzrW
/fQFLDJ8rY3ovpKOrnQu+bH5iMjVxRnJMUydXfNGDBEaYu+F4M1TeB9/+xG/Ot26fZz83RxbwAxx
9+WSyGGfKOEBYNfMOIY0q9t4nTwVWy0dENAs+Xcw420kDN4zVNfSEMTulmAS1Z0SGY2uorEszcKu
jU6AEj3qCnDwTVHLKJc/Y/PpAzchwB2C77N2kygOxTz2RLZRgcyFG0ccGROAc8gTQtYqtqbSh2Zz
SpCNZ9pnQ/HxUn1ZhqXfnrlNHsltcXscL9yCgPR69BEsERuqNOiFgewrdyO9NCqK0sA9HfUOw71H
/0cqm4WueF+nBtLQHP9SeQ4glBrs0/2bn0ogKBgyF/2fqgmZ2QWRqtLjd15dU70ebWiRSs+s1taD
6cylhZNLrgFymiSxekgdSl9MiQulgkyDhGd1G4Fi7Zit7w6M1uRcLk3TZIRRvcVeCpwve33Fc06F
rPr49UMKCJQlVjvkuBRJ7lkc4CU45ypkmGE9ALdVNlcFq59Q2VbmmUWQGylItMdV92+vPv38ut0U
7y5dx3GCPgaBqvOwC6Qpx/ASFjkKfQ7mDw74YeSl4on3eL/hqSqK5rVfkJUKajrVqYB/smjjUS/Q
mubOyQEWlg+TvmJyB/NHz8swcWtB6FhW5OYvSMPSV6Rk8jY96Zl4Xl3Wu6HWYid4QwbQwV+Yfzmu
8wMnZ3XMh6xJhIv0/SzhXVJ8SHu8+9N9nXUoEKfV8q573KkqOkVtKHHMPfvDxTKv+IaSo5Bqv9Gi
YgNXUzJjwJGr/8Ch+VKVLvahGM9Qz4JQ5l+Zo1qSGndY1i9E/S0Ac+mZEk1woZ1qiqtIAMMR90B2
D20a20D3qq7TUYEu8udPLJSR1gxbpQuJIsF+pA14g8NCGq2OQQnKVisrQ27Urf72q4nkuoeyINzx
i/c/OCTnfbqVZml7dLI0L6cx7hMGxDqxKoN8ouk+EtmHiDdO9qwDF4CqXhBfRac4Qcyc7vY37AhI
CWauYvBxs9Ji4/BIEPl6RZL0uOxs1UIX907u7y/d0tqIUoTAl3P2sBwF9B2Md1gztC3o/dviNm5/
Nqyt+7WyNGeRcdtGu0ujEizb8zoHl2GAzk5GlCzpcTZGo4QllHbK1nVjOz0Q/znfPkGTCiC6YpAZ
N2npL+KAt3PO2Wn601OudFUovw/6W/5+EKzj/urjfP+zI0DeaJhGyuZyZqVPYmUF144+YQAzOCJA
mx9X0bjbnk8F00b6TzDCxozCVxUgQrOnllk066FN13K1OXRalehtu8NJMgVNWyN9p0WPwo6tlI/G
BbgHKm/XBIcgommTMzhTKIqUvkfWJeE2FDtm+MBXnGMSKSkVreuDntPI5+J6PAsi22k1YBOplPVS
IZCSY1z7Gz1FgHvcI/XQKRrjbtke/iy/xntgyeFYxRQs4pRgDM03/QHBh/l8CRtl0OK/iTfp/1Z5
7HaasugHw4BOi42xdA/quYFamtAwxZeBPj98cUUkc213T6+jMJDm+Fko2ja1TT4bt49OxWo0SA2e
yA25lwv61Uyvt1DyFumeW3rcDQ/JcOu3G4xNwCIxbYCiXLR0acrL9rOUBUt4rUR/DRByGjIoJh8g
Mm7z5gYjdtmgpHVyUceh/+AXQQHMqVqks2wpFI39pim7Oc5lDlN08scncOzjBchUMkCwZkTdL3RA
bg6/RyNpnwx+VgxKGj/sDPg9tEzE1W1Ieoz05OT29CL4g3n/viTCkNkD2pHsYKOQrfrjlnRpcAln
dtIkqqQ+sHmcn7/QX36/9GMCV03/w2oD3it0RD8gudXSmN76erJzpzpXj3ybu7a+oCeE+oxL8KBb
yz+hFsuGxy3uhGZ8PRzExg9xDGiT5P78AzKmA8BEJFNQv1sMHdtWaSwOh3NB6/LWwjv+LZqezzCg
Oyv9KAwU5fgu/xA0b7HqxYmD4uuIQOaiNX25JVzlapr5RptCoDO0jdzAIyZ30YwXJW2ka++ZuNI9
T8ZPMsThrPT6qip8iAH9FICxXi8ixW3bBlcPb2IR87dM7pCnzvATpqeUxwPEg4tHYZbNTF8CzRZR
5RavOGJdiMW8Y3qaK7D8V8PsgKGgiilrQwnqO1a0DFweC72xm4rnk4iBE2vAFTyvRVT9Lc0xDI4M
1M4QydaiLbzIQtEqNcibUCaowXeYKjZU4uWfww4/DL+JCGS6TL3L2ofl9h3cFE3hE0Ua0YiNnJdK
xrn9+QNlWmyKCrYBM0lHj9MeRNeVm2EXRIqmOCBIRS+b89Sxc0SsYmu7UyQQBPb062SIEqDn1YbJ
m5VkTeGDBgp89LOGmCfpVtT+4ngoH/BF9VK81TNRAdE4MpkA0H05jjMvr23b7BPicp9qWJyD0C8O
9eEphJ4P0wAo8aWd2PHfsC0R6+I48en6ZIJNIF8VivT05/LjkzWOl0J3c/+lknVhE8N6q7LtkkEw
bwOHG/juoV9sVfXNVWDBlnYUYsrMAtMT0snh9+bRgqe5QtQozpNPOz2ZVjVtkcd7oObJdadTYVKp
UoSw+k3Ya6509elf/gZHIl3Qgaw7F/Djc9LUAM10iju/UAdXC1b8SV9R8LreObclyMURZUwpXQ6F
jjP6xAUFvHvbn1M/DpKxnJvMxH+BE56wU0WiXZ6bXC0okGGEDB4RfP/jVcLr8Ev3Z0ps83e9Vq7E
i4BnI91FuxT7MCcn3tbeXXZLGShemhZaQVw+zLtKfjz7ILDbhon+/B6DCEySKoaGV6nPeK8zHAof
5bebe5yQNlFrqZWB7xouI/lkVAsO3y0LfyxzWisKOGmi6alQYHcJam4nY+hwgFiPacMZfR3lm/zi
BkZflnOs+FxDZhdYscOGpIh2FrCUpFRvTxivcyrXXt22il0jPHUlMXTyE2lc+hlp3wN5A2mPoQqb
BLsLliD7SLZXd6cvsb2w0bnVSsvedirKPQhu/+VnBijLqiamR1+B3WSYfN8w0id/pA+z+RvJDEmC
r6EXzYmLn/z2jQTCx69ZDXIWgoQ6N/nL60L9zE8fMuHpsUO/8iQVy0yAOtKXDFrX7W0mpDnWlH0W
ttL8CeGCQpZVPNvMiL9u4LhQMr6WuacoXbekTADBT7Up6JjAV1JE57bQHtcc3ow5NCSjHh0vCViK
p0Oe+slwZ4lH/NTbQ1xkL265+IGVRjhP04D91HKuL7fcxSEKpAJS9pTIQe33Tad/Hp1bOmxk4/Gm
Wae1FAyM0FAvTnVTZWKiHcStciuXih3Waaax25OMVvjwXs3hYF9TkP+O8YXMcpg8JbYtCRJUFZUf
01e+4fdx+hAGuNbWvR2kgfLDsVYTZjCK4oM01Zm+BMNell5mshM/H4BfyTx+5sdb9ISyug8RAR66
7Ipy88q/raWi5BDw19dBCyn4wk9NeK+f/FHgUZXeg/b+9KeoGKXo24RCL7ZvrAZSKrakMtry82qE
eZTc2Ot0l1ymN00q7NCFq7wHLIxxXNJWcn79OMXBdMCZJf+CoKO4qH3sucxil00jyrCd2h4P4nJP
ak7VwWvtnHO6/hLQ6fRHPxJ8FHSv7Y2ri7DG2pjlaUa9tDwdCSdvkaGU66DxGHjcqxhhYEfkujYs
glI64cRbE/KyVPU1qk6ClDgxZLB4pX80ln7kzreP2Bwat6nstyRYquV964A5ZTp124xPkEGopxhm
Jb5UKRLx72plpuib6kOsbadjZEPdSE+OCucwUSf4SyIYT58PxCNP1P+LCF0Zkel7FtpA+lNVCILQ
jfZxp2a371PwE76Ysq06DqHTGAUkc1nWTp02jEZqWqFxGuqMVM6oSXBwYjXV3Twxx6ZaDc1+1lyB
9UAS0eqN480uNgiK3/XTPoGwsrTpzOLlTRJvhLOGadavrN6XEydQD4QoVcU/CIHX53H+hzfI6RMx
ZhCS08/+3obJfOuxvb5i9MZrMQBrSFVdCVfr2Yf3Vy0sN4o+dEjf/J9tyevgHqZ5eC6lfNrQIqVB
XbKG3lyvQj91FlkBHOqrnEtRaDuslgw8Uh1qlrJcZMPSvihIKuNP1SYKIOPOGhTtjT6X5sTmfDlq
FvQz6eSQ6FJJxfs26owBCD15mLhHu2rwPuZ8PivHuKSefZOAdj4a7mLl5I/g37e+FUafXVYOqGuK
1ZDczVBpdQ6sb80vFRZLPot7Jtv2RAXnfxWIBDhcx1+PiWZ8o6iCvUgIYYVPZPs371rhEGL89Bca
iktDShSECQjb2JtjJ1M/GbcR7fwT6FjzxaJpiGc5THCiWUcd+r6HpDfDR5lVLfx0XSvLrxa+O1Vf
9pw9hwQ7Nd9Fj1M0ynfFOfb4L1siKi2qbUk3wmpz2u9ycfIs8bawNG1GjX7guVT+SI+dzu6AQ3Fe
0Fx3jAdbYWArYaZ3y5whDcMM8JlkegJlEdBGMYEnwjeR9ZkDEoLoCOnoMZl4vtFKdM+nB1XOzyL5
DJnsex5bGeMaA+l8BD8xsShF8qmlnsw3+a3G/c3/tf7dDzfzPAwP4K2tShNkceMiQvN5YLK4pBj1
2lLMEm/+LqRjfA3TPxV3XcSZ/oE7dwWRuOPF991/BwIhzELG/FVj7NXA/u1FyKzrfmF6eoHiORMR
quHUxLk8oR7h1srcH+St7zs+FXXiQe7IwkhDZp5vKEyKehU6dByi09VPMjQZsSdVDtwT0/lEXD16
iulXtPQYEvK4nBCgxXQUWNM0BwREj9vGg7z+WqGS7dT73G4vcSgNAelieGdomg0BEWaK4pHki4t9
fuSWTcyICkDfnGPFbnNB9dFdL8sGoNIGFEYFGNEf7v5R8REn83AvNG6jguaAD7DrvePvLPaTHagf
ScHDr9IzJN/ugVe4FvJluHd1Yz2BYdbO+NlEW0cXo08T9ss86WmacRdSfwaZzt+OL2Bb4wnqFhPa
rneGZ+XerNlT6xLg72mBjl704JOwWxcaHZwoQkN+ZYWyoKgISil49iaBudWT9OrqdjOZMpd+9QrI
uek16IVxkqHGrsDmLgniel97kSAPxNnXWlNrtBB8gkspiPgKSWWW+XgWdCSCcnIL/KtO9fZY5hMV
BW6DmOKP5Jz9a3BqaE+1BZWCT3vKlLsGLwF+pCyuamJwElF3eoGPdVLN2+xxp7s08vXCi3t9YCYg
gBejq0DpOHrh/IGtjasN8FF28z0/9wXMuMnJ4LvY+SnlHpI0pGsNRiYFkIuejYaYioZY1+LhAGfD
Mmy88/+6l90Wp7n60OIuj2HG9uE8WP/JJMkyDzQZUT4PDEVcluA7aqqIMTZlcX25LCf828LXMeZI
VrIr+mb7BNDSeqrLxh75CHkTy788pnQC6btU37c8bFiq9KeaFPPmvgnPNZZe5m/F1NYXds5jLIFP
BsHmPQB17WSKWLXGDIua8senrk9EBTjfRgXA7w/zE9XQgy6kP96BeqweAJa/vxqtGOwo20Rdm3De
hXuSXr9ihyp8gtb76o01Hesg/0VdvUdoJ1Eue09Ta5T2m5Nb3RcqCg36bWH/OHbJoQvRSqnxHU6+
XMxufJGZuDnyVF5M5cGrt0txFptJrNntz+aREXWepJna4osSrqQKXiCCjnb000nfgdHPYuUb360z
E/EGjUchiz7iFXOsdzNR+r3R2slhG2ttcpfte0NNhDHBEIWC0IQ7BESUz43RQk8mc0Onf9uDXW88
Gy2PCWQHBZmvxqBFCpSd8PsLXlpCA4nDM/NCTU5+bR9z4GoFXjw74rlbDfmqPo1jII0xlbaJDDsB
0qZoNMFT18oBqn5Ep9mVhS2s/WktfvscYPEUKuHspvwcr4pnbH2fC93EHMuHSys2N0yjts3txESm
FZ8DzMyYeocCUaxudNqFQZjsXSRHaMInyLJytg84wB5/QcbnUaDWdIjDLDSm1PCOi6rSJJDGEqkF
FB3mJN7SOVnyJjpgrsDHGEcsD2GH1UmX+pjWkxBSYqPjgyk0w2OfGbJkpBDcPsZ2pvRKN/FUkjE2
KR/Az4bDlv9pcmErX557PeMmx3klKuyKmIZD8o6EVR3GCRgsUlLcoZ8AK+MwCs1N5G6hJMxyD83R
uzzq3lHMbxmQ7FpYkQOnZrpdVdRsY4GItMgV/IMlWyCuyhvfe6TAZUacBh79yrOTNy+mDo2ZaTES
xj1EQEUysWKOLKbMiwjS/WLTnUOLfk8ypFkoZXQnFI2ASTTnjeru4q0tx5hMOD0tlpbfF4XzzBP7
CPZv8IbUKuaER2NP7gLz9+3dEh1mMkhxNiqBHxYQubpSsMryfQNanMuvn4JenTcHVBllvB5Y0X1A
NLaF+HK2I/zx5A7Dt96Jzzh4fGfkvWct9HBOvBS3ZYRzEvX9hnt/+S+41asUsG61e6rdHsuhrKW3
YoAKwjnxf1x2ZSjBY27PQrw7OMtmM/x5pmFz6ThDGgDGQ7W1p2QBEQpDYWTxBPiu7PWBy215ea/m
ge5L0Ly0BqFJn4le0TyVIkc6sEstWgNA/P5n4n62XdQxdmEGVQHh+WZFJCSzsRGVvmnPZ8LEq1rY
v4l89NeAcwbu0vddKEw7LrojtFNTgG0hlRWUfEeuLDC+3hXhQVUKHo1gEdPIloan2hSh/jliL84Z
FWPhCZUbd3G4UpP4btb5YYudgfBHkwXWdtsURMdUD6Z3uQVeN3lHuvODfbNqgflbodgnq/dTtGfF
VHPWOS0Y6OpkC45UyeA0KVffRdRhdvMb7dY4sYWrjP7K28RppaYAbt30eeGyFeNQvc0QGLEvI/uD
vkhusRTj5mnNvwz6XkoxO7DKJ43ntM1EsJ7biOvZCm2f1vIVA0urRuJqdS9dxSMQkRPhuKDxLsLy
43RPpNoyJXgl2DK/wh+Sb8Z4kYpepwe3ZtqUpcKtyidh899SCVpEk8C6iq1nuSCcKnqpgp3Y03XE
JhYvpnlcUC8GjZRm0G75KVCqhgyYMmIgupGUhncyTDz3Q5BEiTLOa5a8qXnau7HEj++2zyX3pY5+
yaxUewzXMnNDDERNmussGdpTDYz0bNX3PhhDLxSbs4qRq9SdlccXGBsNMBPPnhXzXh2unorJIplU
tdOlQo3j8jWQjsjSJo7RFN72OWw8dqupKOv30131wJ9F3SOeCZmiRqZBTYzm9frxRPfdITR+yT49
9Hf+Hj4Hw3YgZ9WzClwwz+Pf0Cez6jonjfgRhryUqrlzVNGZEmAtpXqyrikUZj1yAil+X5oPjtNJ
TqSVq17SJlWVCe1fed+25TndXcRVPCZ4/qcFaHPg6mIUSQSWScDQU+kgvDA6/QyXYpNmKxWOZFPc
nSWPd/LzVp7DJtABMvC91LKkpGo9ll09MnyxVHaciTTDNA2jPeI7cnS4YM9CRpOdBmM76QB/sRoL
iy82yFBbEup7BazWqF6jNxTWjRNk7Zt2mxU8fVBonmvrQD9tKZNlrtgIiNVKxvJTk425A6DruFEk
jLJG5h8MisVmjahgszpNoaXAqnaYoHn63aaP9JZ8AMwWjlktneWWY9p9VNr7Nw5gnkAlzfmd9kBa
RIQAb9zDBo+4YuXgr/mrWJ4CkkonKR7EJNnRtncakDMI09NwqfoRk4pIQGylA55JLiCA5Dearyg2
6gqJdQAGWU3TC2HziKqvAzir7Mzh3wU0jEZosmEjyJ1urBLksTOw6+hvDmklavFPLak4LRc5UgPP
3buSgHiF6M+S47gfTMEB6jSiWyY2QDeapgcPJ/IAU4lrw2TmID7OF8twF5YX2E919je1371GukoM
CmgPESYumOwwiiVjx918NchUpjF+t5ckQtt6sUfRKHTpcmdKlGVYoBvX3sjcRFtU8w1rwMPwyM9U
jSuKuwK1m+C/DeTTQP7p3NXyZg0w6Aw6gS8IeX/B4i8LUlIkwuo8fUBw7JG+mhZ5Z6WhytM1fHlh
GI4Zc+D/apGo58hhAv7XY7rolSVexdxW+PoYdRynIUavRkk+sR2VVBzUK+bH23pLOnekmN0x20zx
XmCFfEK2WLLLHgIEVJy1G//IEMeB+h5JWEZ0iTsx8B8pympAA6rbwSdhbZ2oegQDQQE01qqqvvqs
Z6mOCLK/JagvjBo7FLQ61gafzFzmVyJQdTxj8+W197p0gS1fi0kk+9luEKKvt13BNsPQpR2DRd6y
q0crBhSrQSIaKVbuM5PeeAWNBIiV1c+7gXz02gZtslNbxgt0unQwi9xN0iQsR7WVQbPYCLieA4Kv
rTC5DyHbtvRbBJFYmeym+zMNlIWhfIplciryoNbvsiRaKgcmLmquoytvN2S1KU7gq4fYxmutqkI1
ZzoMr0oocv3FrFzkxb8Gq6NYe2fPWAYgnMgwRdB6gSqJx8gUMmEZTlpUYOOghGuOLGEOTzi+OWwD
KAcpsFnnPOG4uw+a5DHwTzSokZoK5X6Hz1I10AdL5XbGrmSa37hwSRLmUwgkTd0E8CBn2VKRUorg
fzVFqopdhFjXi9YeEcEqFnCGArqSTj7OX1WZSjwCwHVmT9os93a/RMqbZl+yO0RWtc3PAizLW5+1
EF8/ebpryVphT6HT9ZWvYQl0QeDIwcbRq9uKpoS1Q5CFO+mA9Pdz35cQkWOgsSNzTieSSGJ9+mfB
rttUfUobK8ixgigRdzgGFGsid4QU7UiK9/fYJRU73Oe7s+4clx0A/Tc/w1jt7/Kpg+VXkXI5/lKO
bxFpWDAblF3baBtVNRNpYTTSIdUiWvvW1WiHoumxd5Zhf6F6ph8+MncnzjApiIT0K95UZHGp3bF5
lrxE2a3Z2tFCWPinlk7q0AXz9XjYGUP+G1RhMJU82eg1KOluKLZTSXKnOuMdEzsyku1mzChvE+t7
HadFl8z6FktgNl0LlQNyZGgqGN8jEZQbWqGRZdLSK7E6Ckyb4xCkEA799eQ7CdYakBwAWate1Uwi
5ngpcfiWqwrX6l71xjT3LYP1cw9IvgVHKzAd7bu0MFLwy87xToBV5fveBmbuy1ZwZf0Lk8kIQj9r
Zd69VnTAZD3gwSAKgnVLeYrJ+AO6ZlRi+Foc2REWGTaihJAEpYPwJssFfuVLsU4wKeqI/t2L0Tu5
c5LXlpQmy7Vj2mbBBO5Z9Y/ZZlYu31HxLwFGdtrf7idv3yUGwVu7dqCxRqNtprwjlEKnTTUmcO7d
j1kBXo8MBk4tzDDyDzHSS3hRdUg7/MCFVArgwjkLkt3a1an9SxCWf4C22VUNvUALSjn8R16lqwYR
Fl3BBNmmuY1L7dHCEFkM5jUSdTctj5BH6j/7SiszTXMrLAr06bC4ONJtt1PqhzyQqzHrFnswIIht
aWbBnxz8zl3cIwzQpSYcAIHhKITX6tPUCFftiduPE3IOfb80gs9BSWbsENCl2hEE1mfPCmE1qczp
pBTsjMJWhtWiJSyku0QT8FDl+5uZUZ3o6F8X25KxF/feqdCqE8RgCLXn0nG0UOXMY7cpLTK7I5dD
LTiy26wCxzlOucmKVaS8pghORWgUkytoQtZJ6uAA4SlEpnBt4VL1iTE8sxXyGrHiQ709Zsa6RYvM
iNxUWqFcnOb+Thf8ifKWJtyO0YYQudxHmbZxNimUp7psyqFO+UGJBDllBXZpcjjFCmMvx9cScmCH
hS4keK5D/vky99Sse7UWP80xSsjL2AT+ngeY6HRcJxvjdG1nwSoM3b9FkcVc3cHU3tiXW/wucAW6
JycztqdpZXVTmOZdjIK7/xf5i/06gtGZsluWC6WrmOGxW0hFNOCD6wdPJCHaaBtHcGAYU9oWvHg8
5buuzlnzxZrJNswwRh2VB8oVetTAyPocXlocxwo50O1OTthCWSRsATrzZs5pBHoKmeQIuIvTZdfw
uZdXxpZv9bCgrwoea8qd0fGgnTX57WwpFoihoVPUK4/trM5C1dnTUgcw2wLSjlZLJPCmgoRZWa89
2RYhwliKlvfy5bcVhmFWMHPGJ0vz+96iqpp97YXbYNlUrVU2gn/vy13UwpDTkc2q0GF8upBE1hWn
yODbNvjBzFD5aLFeGvP+vVu1Nd47cDzJMCF6xY39fWJOTxvekFCO9Enhqbtx9yRrwlHS2qa3bsvq
kBK9si6O/7ZJVFM1fwxP8IBX8nuy1LzeivbS/wTLNnmCjUEtMklRmg6tRDYpjajKCCIniUC5RCwu
GnBq0k8PW+9zLAiRxASyiIydByJkoZcymB1A0qQXLDHUpAQa1lL+X90kRA3wYJWlDnnuziR/XFHa
hmlQo2HA776xxQkU4Rn1Yx6f/lUgdMoWtQkJDH4HpyuUeR0XrQPY4nTfAjzHajehc5eIlx3kdFaL
7QyRtqfoOv+y6G1ASklWI0nGqbWYnq1qGLrvaIRo2Up1IL017au8amMhfWNbazRFEoI632PUYsxl
MPdOjnImu11znleI3p1sTRjT0rC6gFWFuMH3C+VT9kTy7OB9ZBf7jpcpr6t5WjRHjQzgDjqVNhIX
J91pMwdBlP4V5W87EgLQ6yYRj26/4tdu65eoLe1NhSE1y4im7y4zMPZ1HkdlpWbuA8IS9ZPbyB1P
zfoeENdiDvRdDskUMjc/xdyUqqHyQ4DzITLg0d/tAvrUHvZ63Rlurm8JDLCYjFW898hzbXyJYH4x
QeEMSNptY/OiJJ0b3WRAy6EAC7Ttlm9jqOsPF6dzFPDn67D0yWGr7eD/rQJ3lu92zR4u635za4q6
8ufBNgx+o80Lm7A6dFJ97/jPssuQsN73PO5U4mB2UVphEBQaUiZodSzId83gGMGZ4BI6APtiqFXF
uX1EGz5riFuRCFQiIZHA0wU/gMt5gJConKLWbSx5cenL/ve+9ZV/eDBZ9KSVf2gri8usH60CGPuZ
gPin3M/Kqv/0Xj24Lv1x2eMF6KtnFHOjP2pYLl6646/gEXpT8Y7x0zXb+E9yDLXTuEn2Z7BlWZUF
GfMOUftork0b72nPdEBk7MRQsM9Ny93RFj/wxxfZLDzNyiQrIA0a/NwJs5i/24KhOlsuKOy21w9j
d0HAEt6amqFpDadbRNiDgsoPVWpuE7McO5mVxxPLtAIjs3kuhNPw5RM0JtM6FMlr2uDMgkWyrLSp
bBjPLwZ+xKRXJcktWVn51tI+RELhXdefMoaxCJ4fPa8EsGeez8zLmMenO6sQtQjfLGaaymxpur1Y
I6Ub7NByahiHGFo2mFW6FQ8DbS+4oLOT7+7EuoyqvCzKvBV9lWDj1TXfbzsv/8CEPyyjtbX1OEM1
A2ygctrYzDu1QutPiTxJm+tYfllkjWByD4/o/W5RTpOil4Kw6+LsXsyVyne4XhMprzOeOnuxDSIG
V8egowoKDtZiB0TY+LCvyKIOh/11W5ZKPwsHsKtgq3nb6pU9Wjw8cs+S/JWbikM/1Zcly7mDHx1i
xA+LpbuMf2KW9p4w0zPpceZrPVVJcUowpudU04hfRYPIZYx4+NVxB3w4BMduyNprbefug0+e4WeN
cWMilLN9VpyZPlR9BeidGxYCArm2E4p29d1vR6OVcdatAcKpBISDVW8ecy7Hdmm8NGiJUpg2NvdL
bB8oeX4copyi0N4+ms7saZduzns1rt1bnXvv7a7VDExPp26LxNGRqbnpA9OVTNXVBKnRBjILhKa5
Og127Y7wgo+uhtQU+PIHkcG5hVbI8+6UONNkqVCndEEgrchiPqExuzmZXtdFu57XuRnoKAG0raUT
GkISXz8AN086V/7xY33gJRBytdkz7Nc/euG9ryBUIV85qKdD/kQEDa4RgMeiTDsKFXTZK/T33WMT
S6qCOSY2a5EsuEjRv+kr3plaK5yg+O0dYLXBWWSh3NP0qm0aqOGlfSCJlHWDGnGspg9N2SGAEKwY
yvY188E/uzTE4i7eHtZ4mwVcAfF3lR6amDLpnbzqXQ8IspktJ6eXkmGEIstyYzT/cTXyHF4K3FRb
TW+Rtofd+j+prHhoQdMCK0YZaGLPyI0LY9pWdjlZBTO4s+lV0o+Jk5F1jgfzxIjVatSCIVrwJEjS
z+mV2sbQV0QkVb9wYxstb6tGeCOLDPqDMwNcXFREArmhUL44o1NWXlZ9v4QXRanqy9V3bh9Xid09
kQiP9abq7YnDTHHy1z72jPAdTjjGPz5Ww0xWy/bYPQPtECZkz7n2VTNaKsLqXs4pR94EQTfUeWf4
Fm+2kOL4Me9cbhA4OuXeZS02Gt6vSZvXo64O3tUtWLIn84+smKwJ1/OeRkAyH6VCXBwIiuhSNgdq
r5sP8kh48Ltm7IU8t3neKpdEub0kv4W6MhMLVcU1Wyp+cNpVp1QBG5LzPtCLaVuR0yisOa3TGd6u
D76DscdQZ4qAznZKKpDg18um50/PpEZt6zNbXVoVUiA+ioOpUSNdR5ytqlUlTTkeoOZoJRCzko0z
asIuaJqFJyAm047Vhom0f58zODn/TzghgJU2yN5LpQ84NN+sRjR0EeoU/2uwHtqvjeINNGIxTMLO
wHB+QS5dkaMDypGvOLl5HXAZ6joj9gLmuwUN/kdOJuoW/uy40bIMsnllmfvN2sGYdCFs2vreY4Vw
UyETAItWgudOU1F7MLtYcsUbCRhgHecKwxcTaB0IWrGoTJxWS6xeAP1KkPgWJWYTAnhcDSremM3Y
vl8UrWhjcEoDYj/o4tlFeONhsfoQkaz2+OsSuwELVlbfoLBk9nxgIqGDFD3WFZBsEvzG8+fDRIUg
bcnOIDTf7DI0wfq+OBn7R3P2glYMX7NJs5N3oema4h6xz1kcnop7B0AR9ABYE3DqlJa4U13u7R6e
9ev2383N3eEWPfXJVqWzmGoGCouZOdg3f6DiuQNDsGzjxEWoXjnYMQF8kqfDVQ0ndBjKK3Ervkmr
rVfM5ZKHc0dur7pZW5+8eqscHN9KzxBzkx+qp9giZpnYWwRryvGKhXqKWrNfey58iMFAWfZ0xV2p
g0LUErzr2yCkMsmsd+YZGJchhCwjQ9BKEd8pL8z+yVWXJ9wfm0/Fm5IBYSboo7KiJVq6Iz3yfCGa
yleCIejq+0FZUWo2tX87JMdAaKKqwbnL0XkET4ZbAhLCjgjIX1B0UwsBYaNbEuYgyrcizH5zRsPD
Jd+DQ1p4jJRVMD/A9MiZrmbjz/gbJafja2V/RAkRvzBU2ZrptkxBbVyNgQq48CDeThoZwi6uucZ9
OL9ney+K5wsSmT43lFBQlOb9kzlkW/xeDDuQ5DiiWCWm006KJkkB6h4h1C8P9n9dY82mOtgXdnWC
bHrhL4whuMuQhwOSTHH1iBwe1UvO5pD/mFf9ec7y8RXQS4QglLLq2/oPNPV9x+sncjKgxW2LlDb9
AT9RpBQrDHkXv7ZGbdAlVFhEfBug353xyVGos5cLfn2XtVRE4DBcxiRAIJQrtY3BsWyk/gZTWTDC
bC80kktdQPiAWFh9OknA5l/ze+wT5jpNYQyo1+jnzgh/pHbgbbRJz3J3AY9Xzv9WRNyabs1wQxaT
C5Jk55ZnR7RxDljk4e3JTW5tF/XggCOXRGadV3j0EWc69pIFqdOQxbffr+5m/U1zdVi/YEfvVT2K
TjdEUzPO0rHWoSK8rvp4oRnQf2ZXJHygfBUw19SNeON+BgiCfue7+wF5iYHLoJAUhN5tnxz4hPsf
v/0XWJ0EHlJu5GkC/QgwdQdgyVZaunNpMkDBw+cCKHXR5suW1LbPCVrDA9HlkPLAw3wSNbv4+njS
HQf0MpzhiYVFeY0notrtulwk6K7GK801Wky/vtjN3T3lPP/wRO09XSK85vzxsbtZGzct+gPd7KdO
F1nLaA+neP0cs1g+/w8UQBsB5OaeCB88CwaApHpz7mBNGz15WDbNL0IusHNVO8m+93MmeOVLrpeR
ymjCUHpl3tUa4sSNWY8DHwEZmcshuuVskcQINcQLIXS5/GCtqRyyhKMNNykI/SVRK2SZ5TxiHgqQ
DM7xG64vCMwuy9/pLhrbc+afe/Pkqqnko4chg3hO3ir4yYCYLstWSaCrGY+dd0Q5E2Zs8ruz2Cxi
A+N/7iCCPqvi+KoaBfynH4ajEgsnBOshu1NHx1/micflB1r4dnyF8xRYiy8/SJ/sU6K9hgVnpUaQ
vSecbx2dzKsyIGD6j+HbUlTspoRs/qamJaIuCkezSNQJoacYLO/cjjxlHbz9Tu5eYjt9CRrh3UeK
9Wm3GCh8Fsh+wfY4htHLERPyiTUbxKGLQ46fFtPZuRJcHRs5aonn1PdWDcmNlh/KyJdWlFg2ylm7
xJ0d+SngWMkG+GxLgrKv4J05VwPExBIkkbE3x1KeCsTL7lUPzOniTwy1ww90LK0rJt+PGJQwIBMo
61o815x6Llbgge0A8GS2rqEZp0GwdmLnF5oTWhjFr48XHOmFfLkJq69iVpGZomoU99s8ka6CmDcj
vv8DAKIWGDqorhpZa+/hREP8Cjp/u/qS9gt4cyZP6/9IVlgFUFnZhHhOnqWasKc/PXXLuYsUgKep
FLTPJjFcj5h6fy5DaWxDGfUPJRac4ENcta4+F3PChJ5CZaj8xQrfqmD2ZA7YQHCS9/RB8UnzAv2I
RvjoDyOHNmZZMbFKzeOXnwPY1lmOMS/TknVGc1rB6OrPYkN+SMKslGW7iYCETlahuCYlhU3OL77r
TYp/731a6o5oXFhiNdCLQf8NvebNiMS+Fxdwoc6b7gLgXuNjQXXCWzjKubpOfsVCuiuNPKLo62S5
9afM0kcl5AyIMwbgwNRSoD587GAKqONQaG0V5MuM+FH7KbmX3k61UE+zpqoS9AztZKq8xvOAlxGh
PqsyDRskKs/t20iHvdoYr6f+C40EsTpt0IYXB0KN1t6fM9ydr67GBg54sVwNHmXSeG5pfuRygj3s
9ARq/bUGlUhKNxCoFzhEmaLG6hyBkhMJatK9zGrGRjKn4slPdYgOXV0rMLPili/iFgA58sYlc7PW
ji7Yt+O5o2r6Jy7FAVndu/9MJ/HQBdhXoGWRpFvS0VJBR+Zv68/IkMbe9gvi+rtz+JfYkZJj/VPh
P9NWn7osbzJuzokbgnyjuHJCCblNdUvro9Ive88u/aUiq1E9hCIbOTbXe+ogKi286iRo78Lmksv6
qZdWWO+upsI+SGe1se2IPbMu/J4jz+I1rMr6BISiUBlOQY09MOsXzv/Uf5dGML+kbA4/uGxVXkgn
G+lh/fuY4hqIwbLGEr2BYObtltyPAamIMOck14nJL5Nw68Om2mllk9nycnghMfy9vEUR+LGz8IxG
WEHwZPnw8OmZuuJ6wPHhYua9j6v1Qu1yOK+VnNBcIib9W/Bq+XijtmG2xBQzk+JKGMB6o2UMQ0zP
v/HezaokXTdZhTYyPA0Q/jDeiumXKtkfy2hNoS6ykH/DfzP7zyXIrP1q/UUHRRt7GPNcbFkCkA9j
7E/4o4aejnx/w6sYoY470gupeCqn8guP9FFVgTm/vuPoMlYHxNzz3UaMXYy7I6mydgDwFLob6xVQ
qAGpMMIfbSpU1YRq7SLbL0ZcxQgbenCr3jAjZBGyqmEPnF3Hnmu69ieane9QMLn9kQouMeJv8W/F
ULO++v7Y5XrCbf7cbhtBfy4BuKERwILs4EOI+GACpthsHDRGqubsC1QJfx7gHZ/zd1+myPJoUAZs
ECSdPHrblebNnkzB9Kxa3s3eGhaxjzUV/2WL4yQIvUJCGP+ufrlIR1Uqpl16JYgIDcJWtEs+JjLF
/uhDiHH3mU/Vscc3PZlfoZQ9jH5gAuWu+9NKdco6vOdtI9zUs4jhUmGkkRyp6Bm9QiZeNCO0rwZ/
++68YRb1J6oRZ1X7DaP3RdjgeXIyJtzrDlCUFWI0CsEFpH98P8hdJ0E2380d2+xKtOoFnLoPymBX
ogkdgjP3uv8RpvfreiL0dvyARbFXNAr+t/JQoLSYVFY5YzuaAos+Xgvf33iJKpS9n/dBCJwhSAZS
E4NvHQhNs0jogWwkqGQkUqwZz95ooHjdEFEwQC9HnaihJTUm2aQNVuasM2T1s3DHPPfvXJdM8ICr
Y2Xlm0JSHRayso5xPaRCnnTb9sAf49IJxhXGkr0YePIpeKOGjTyvC9WKkpduHVapat7Wh9yQFU7Q
xCI3WzDnHS7zP5WV9vz7z0evzUYzq7JvNsH3GmaZez17MkKnIJFbVhRqJedz+TgB+WyrSekiRVwo
nAfX64twODj0O4j0P/xe3s5Wri0LpUZY3Ynx/VHuYYAs43HAUtSDDb3n5ZlNOyDuLHlUN68xKpAS
7/TOGAOWTS9PqBsj0sI0kTrhnBXcew/iNcxOfDla1EcIGfqSSwDNgEQhFgG/AxhY5Rva3WwmT52z
J5312tsKz7rJdsM8JhDZUMpI78dWNWjk+rQF2EbIqq3xUkAi1Z5ma/xlTx2pxGkfsdd/ru6/38NY
CeK/6Bu8F5jnN8y4IkxzOF/FhvTpQEtlhC5ev8ZgBJvstsMAUEJem9Sg26nJANV5AGG9chgzDIS6
XlfoONPJCYUC4al/LOj0U31uBiJpfxXCo3S7V4rZReOBiVr/qyUJsMQnqXcvsj8xTY0y3JIoKYHp
U3vf/XWmNy4Zd2nQ3AFRdAZxTasVJb+w4m1CNvHNDZOCiwutQRTlEX4sYQ/lk5xus5faLCkTEWDk
69wyMxCvv+FrIB37wspaZzUJYZD7YQI2/ha0yelSuOvCCl60CQ26IvvHqKuZHm1Wj6bMD2lYygcj
xYVef9fH/HEnD43KGrrUSioV5C8FYhJ6wFGVh/ROPhmEUCq2IhwoZrfVK1DTWkyv46Ntswb8VGLj
G3z3Lw/XvCjQNs+Ql3ISR6CgdMyqMsXbFX62FnJ/c9Vnu1AXa8eKgO+RYWSjbLGRsgC4dxgjReQ1
XPh7ULlK1aFg9SFQTYfDqFiQid9JxGjTYeQM7xnxkGxny1WLHXirJk9d4hV+FxvpzYvEns7CLs6A
AYL9egclGNLLe7OWYT+JdPKeEKEvBMLF1RBZNEsc8sx0V+uC0gK4Tq0CEHkSVvPLFpPY/ijgQ2re
T1BMOggQMzEpKccntb1AFrFgWX/AUjbhs/A0zb4WQIp7mRRHJ6G+bG3rNHtAQpTp3r6RA5g0jGuE
bMoUyM9nV0mK7g7sefX7oxKqCdzC07kkiZEbhZo2u9chqxXDl/jKB7DoUzrrCd8JIDbPDwvWKVak
msU2WTVe6xWYg/pHRqpLjb3QeqwZRZByXoKyhgTt5cKcRwhcPEewGxaZPax40gLVZsQo8i2K314H
Ehh3nFCi/IkbYSI2Q5NnJJw1yG/mCVK/1ImjxKvk0jzQMeLBOoyBhcoL5BD2FCO3+tfFo10xsJN7
jKPlUJWJmqaSo5qAJAM0F8Lcgrp1W1cpAIc0pDBF3uizKnh7CKd5dri7inSfBOaAGCZ+FLreARQT
MIdwP7XwclBtBXw/kYRYXHdZGwOlYSP01OYWZguBI4WmqMKSkmy64St2fwGyU8Pi5FL9yZ2LajE1
bEEOyy2aUx3GNNpNym91/972g9vj3oHMnGOnNm27dFZmItal1HswLRHU2IOa63oO9foCNZydbqU7
ZSqZBBol2WaU5lA8+AqVq6krGfHh67TYLIhAiac4obk7OmicwWHJd35mxhOPLgdfYJdWAjUt+05t
N2KVLDpUa8EzlV//NFK5KR6iIOaA6i8vEoDQ1AUh8D/D7DC9r+EKkCdQnmi4z2xGSzGLlvhXy8J4
UYsS6iwTNbRKABwIWoJQTUEYVu9qpzrTD1HwTji1aW2k1oIFNNuWGz5XujbqodZUgnNNidRHoJ68
RIO1zB7KnpHNNPzyhzwIjHz9hnK/RIRiv9dQtCXC0hndHB5gs5VkuxjPPyz5EXiWTAhWj5T7zOfC
IovmKDikzPBHD8soh5E6qTAxGQ475HgE8A8uke/SiYCuJ24Bt//9EK2hX1wAhWUb4Z/sD81sc19j
bib70ONNfaxesI1hFaRI1dZyxZypYAWnPlJBPjxAzlXWZkP3IQfGBGRIyKZksWh9/FwgZ/EoMkAl
mDzCTrgDF57cVVHYUhE7wCCNz+VV5/8ejP5oph38Fj99fbCB7EewSN//oYUG2Vc/DKRR+FbgTKOO
uJkip0atk07D/57e3G4Pq6rbhWZv7NsALUHssM/G+8wQUil3ii14+h02mc6B3ZiVEvlfSbgZ1n3J
O/A9QtjvU3NZHO4G4wBydboAWCDaB0/JgoFM987OjefB2WHNsvemd2QxQRlDTXjoqqFJX/kfIn20
3IY2VQdixJlXAORtn4AIVa+4JFPHbcVxTryM74ytwtcFzbr134oj/LLdFqjqasvzgkTiUrrd0LJW
A3YYSd/bgVWfFKHTFMH4U801MxKd90nf08nr58lTT8/Gg49TF9Z9d0IekrMaSgJnG6nN4r0cGEeB
4NFiw8YEGnW3LGJtBYzFRO1UcgoHAPXchPC/kjE9cQ1A3EwPIdFvdUhlPqfsEtcnFQLQ/HNghKxI
8VR9ecoOVpEJt1ngCVKw+fd+wKkcm4wTru+N8jb4XQKiFYRWIqZl77OyisM2Tgpi05NwTFs9VxvO
GWOby0jNwhBKBN6o+B8ekmupcM5NZatXkf0BYRA7uPt1qnV46qMXmU1yxvgtaoAFCn9FhXgi0eMC
Uly3KVMih7QXrLSoAPUl7R/WcGEFeNCG1WIO4GQVhepvERff4rxzZX8TKJISP6IRELc5oBjYzfdC
ct5bTpXBvCXMPaD3tsmPYLEaEyfExZR9O3DxxFZ4uSFsuwiRyxOxdQiOSIpqtIAMkPCqjIlRdGty
+icFfIorL+Lx8+0FnBKpcFWExa9X0cfXLHlNlvyoI7wCppyJSsavx/xcV5btEpuZXG77nCB7InMn
tsRcNyR91hHDg+AGrdp5vbZs4d1xmBSofyjHnbVL0ik3kO0naq5P1Lw+kw5LhcSoiexKvIWCCorc
IOrvAJwA3mU7E6BstxJNUxftSu/PTntGrpy4/R6+jaGmi2NSUNXtbUTKgNJ0HVGzNBt9PWkMcqJ6
1qw6/zlxr7gRrmgGdvLIwiwBPAXsCSq+EeuT7EpBCx31R/twtARMoJFPInvuVmnAAb5MPiONTPxT
cfCYVY6qJmYqwI/OVyItnnpDkOLr4VTcMbDqBlhBm4LVUyS8+CcIazk03JOIk9xAUIf+HI04ba9C
nCtWdLdesIeiwWEq2jZ8C4+z0RpYb05DdYD2dUltXwtW/SiYmjpvVpB2LWc4FtaCS9DeCqxcL5Km
uqf7E077tF5hdi85CQVyw44PJQEseu+L02e/sj5i4PaY4msihTrwFFCTO/ma7BKW19VnWPz7+S0T
jODC82dfTHQzDVc70JaYserm+YY+q58sfSaZfCFDfSri8FIsnsS3ti6dFT5ls5IzCV0vBfoaELpT
HQkymU0+5gR37RZdLfSum83t9Kfcc6ZXiXP7hZxk6yFKd+5UoJ857hX54yaHUQy4mnw+n/9wkUIn
lpYU+D2jLr6R9Y73/P0LFtCVPCNzGTt9ef2TT2R8+z1EoylERXlJJMLjZleMgn8/OnbV5SqdgpjY
GtbIRLpZXoZzoCIXj/ox7uIHw9Nw5w7OXreEWyV9bMrWGjxqfX2+0eGS22f+/GtiIxXhn6PlCjOK
p4Opx+n4CgCLjoQko6dJmOVZhxjraRBovTunFAtxFjLceSz+ETRGU+Zzt39kRm8Nk1obIhrjZzbT
L6RCO1b+kmRk1ZCjTqFlRTpphJmEa9zdBt/JF6wZm8rhrLXPozZOV4kIQ2uEYiy2qRuFw4jPM3w/
TG19NeI3edE6jUUFzKvSfiBxKtMGTt00VsZa6jL1x+tRlzh68dS4HIrTyfYES7vOvWW3aLaNM0QG
gDNskYd6yLaFOaCbSFlwPK13taIbNeJNxz7c3tvQ7gYYGmaQ6jH/yu5OEO2GcaSUSrBcN1J4x51Q
37mc5VXtlBLVfwiapMvfTdwLjWZVMdw63qNGhBcr62nR4A28j2ipoFwqp3e5EPEc1TTPpYcqixPV
iOALeMrPQ2rTI4ZHUU8cRJO6a1lDUGHtTj2upJF5/D4IkUoibkxy03utFI8UuxuPVQ9xUtZrtUQO
U7AqGbzKppB+AQbXpTuVT0ttrbi298NXGrkSUxKjjePsphZ0FbtAskwLyF92iGNq5SxTCKQAF4Df
yBxRGn/eJeMYSjxpfvA+FJUtSxuQ+TsLlLrIDfvShKlasHEnPUeb+g0HGm+jOPIvpCJyL8QzDhV2
EnRir+nLBAUrOMFXa8pnVyIXnIWjDXovxlrVqauIgcFbVq6d1uDH4KR275z7Nn5zIwGqQjIj5jUO
inVUDEtZTEufsFpK91ZOddkJLga5kHNZaVenzUiz7LErdhPKK43aT0Jquyw52PzPj0iH1CXiq9nq
zQfAHNpTf5273SDvfNN8jTA2jf+dOHg3u1xtCy8hffkDSwn0m84u0o+xfPFTUarXOgJN29v7OQn9
DuMw7Q42WNzifcUTS4E414Td7eBMAPXXTPxjkfYYNP44FUnZ5opx1K+hN+Sq2XPbEvWLgqMY5zMq
+eWsr//4/14BQRDmbFhxsCCL0w2x9W6P9MuVZgKvV9oAMrm0Ufz/xOGKxJyswQnCnWb5Ie3chNt6
TatTw0kcyjyl47RiVUNuIliudItl+bu/RbJf8fEUYkCxMpiZueW+6ZBx+d7jEQcVJBUTy074gqyV
s6AZ1KQgC3Uae8IUa0JDKhYfj5PdLmwYUwMZA8NOTfo0MWK263rxj8ISuWI9f9oeD5Q0nc1V5yBw
tpfGQ9oMwTxZLebVwRp1mLwql2i5k5cvvQwSOUepEr6blIS4SpHEEJFqR8klrUqgPWMsZzsja27b
TucgicEC5M9c8SORSnmBJGbwqvTK1g4yP3nxfznyCHA0suNTRoL2oJHki9OfUDFb1jVsP7toznVP
tkRjP3yzYCXOCHFZQKa0waMd641b/ToDedjsRHuXCjvXclgDFFw6UDnqvLYLBuU6+EXJ+raa+uct
KUdL/UUK8DvRA2eknQzz/CFM4eyzpJkrJN7InQVuQXyANJLd/UGUFHa7mSUA2OaS2HKmiRNY2C2C
A85TlJq4nBrNZaggV3vrNOJVd36oB82LdHYQpZXl2ojzwk2bQU/zMkzUZtgM19E3rrslFZViBZHm
Hy9ay3bF2tIHvDcK1BgFRvHx1p3PK3/zJjFy765FEcxa0NPsa+lukuK7f6RvgWIiGiRnSgn/j4de
pQmKW/3bmuKmpVvcqpqddq8hPUe6wgk/npsOLXV1YOGGvJyZGeqlsvMqg9R+UzgxSBqT0ESHP9Lo
/NXbd16voWfacXy58CN37ki8Zw1nwBS6p87+XBhPXoSsqKciX9t4MjjwCo8efydROybO/R9cJnnO
kAGcr70MvrafkRIgCamuMEecaRIxA07fbcr0XOP5rTTFVNK2OehX1vdrFhKdgaZHrJocyS/Gx3zW
cDYSXK1yJ14m222Iwcur1kTVnQP8sJkjP0E7vxosoQbGyWwXj6PQ+qD4Mx5OeP9KjSl9uORHaj50
bmVLDqOehW56/x1GX1hnKy6ZgfPOS0b3qoXyQCgEVOeMzkmIUqSX1gIwD2zb/OeZo6XSJ6gZY6yX
HfmARVX8p/AUNbX4KKf14Onnev581w660fjv5KS6DDEjy3ss3T2cG8pTLqjaQWA4ArQQs+BLVu0+
4ZkYk3uWQ0GGWvlyxbIttlVlAW2nVo7pUOYmIhiiDDsoE3PeKKQxpoZLJ7NKqvgU5y7ZI2qosOq7
vMLrTnp2BQFNYaGV0PzuOD7P/bcPYe1wkI70QL5JKnErJra5TCIZpI1i/enPeRUr+uoyhiI26268
zzbubOinXUz0fwASGxp9b6IbvCw5lp5T90IwfW5cGijFJLvdOy9FcU6JaRzXsF/uv2NPwY/5G/Bg
ci29Fbd6dEEdYcpt2xX2O4GT7YZNJ+ijV98AH1ItTp85DwSYSinF7n/OILYTEBh3/5aOlEpT+8An
O406JFdfJ4B2dJEBFMSvDwKgChdXFLH6OLuGqEG/CZn4917fSb5JPM6rxYMnaqHj83V+VhAUDcJq
ON7UP7tPtaPKPuM5Viw8GA+b5jLnIPBXARM74Qva6TgBc/t6emDve3CC7wv/LGZtHiBG6BtdX2Tr
J/bN9ngWXxWkXaPjkwak7dtKCs14LtqZOwzt+QFT5/dWxB0I92XprGE8IpHV7VyAYLH7s463hsIu
rLnf3ZjQ1xaC0NhwqXrgRgPAiUJmprIBORvixTUxIbIZzbhHg8/5Sm/sCsAdsG+rKunXAXM1jfN5
J1W8tQDD4j59GEvO1teqvPyf7t9xXBGEygQGe/ifRYujlqVCfNigaKVUfls/ITN46mmDbsxWDqRP
rz0zWMkB8aVwCTRTyWUYbcawPDoxFInwL+GC4mqIMQ5jPt7Z6hycg36wurBjJcovAiifOyFQGPeH
Us8o5SQj9nr0xI34Imwv9f4tFfDDzJGFejsxOCG+11N7afCcTlqNMGzBda+dAfMi0FipGr/voRUt
DotDyB1cI4vkyxvTR2HHB3QpgswUBLNLqkjU445cDWhTeJkso7g8jR7QG6R4cXB7ZOZ+tWqnj1ZY
eAB/ZxsDyPQL5mpShFzQVt0gqFaXGeHvbyGTwOFCG2kuVTqjhMgiZDk1JYRDmWoo96IOqjcxBliV
FwvlBTwstqO3jMKW9bed+kfkuqXAuES2Id5Z5dj+PkPdDReLz3yDmztTZhMgbtO24ro0868RVIXO
/DwBIBvzQ1bm+CrOBj/KriY16jqIrkH38hgYqRqmHp6ewibnnyzfUerU9fN0JPd6tk3kapjmsnqY
tBGmq6DJiUdd6DgzBGPiUYm/jRCzKRpLxBr695J3YjgCJXKnvP3PWlbDrMdnSBddTh8o9XvHtMoH
j7X6YsIs9TdfPdQuB19xrHrUkxCYs/XFuWeDX4NRnKXC35OfdaAzO8X0oVVcm6MsKBTcjt5IDI4B
gS8y4SFjfM5dnBuRfJNAwthEAIeJ1vwzaCu26czD62cy/+oR3vy9I1Cgo78jq66CUUUliiRCK2x5
7sQEClfPWqJL4BSosQvIA0eg9998kk+1CDmQ+FarZlCyM9aReuEcNpNcxtKuy6t7WTANlQe3cG6i
+T6TThN7RPmd06kJLfZCJ0FvW+jhyEYkmyV1m+ZnMFgObC1yJsZrIRsbpKBIrr+xWm6/iUE2l/AV
SUfIDmicn+77S6kE5bHoVCHLIXgKqmSpwOwZwTItrGX97Uh3Dv/ukDtX/qT5zkA719uTcCFjK+Dz
YIHQ85RMDmKuJAdEUYjGx/sRZ3THEu8EE6RJLZUzUT5SS70QVVy/UHFKsqu1dbTa3ZAAoGS0JShc
u/ZsgZKGNoZQQhadY58z+3yYq1yJH91xNxc0WmZt5+5eQ+dDSnK7tni1DTcluvp3h96FauAaS3nn
JQDvsJyVwAOO5+7cidyAf9aPy3lyuZMgEV5yI7cbzUAWowv9up3wrw5tKBW7K9N00IwQr/K0bK/v
oeE0ku9Zg2kwzG2XUN4AeBd99fcfYlVijK86Q5VsQM2LcgjJAH+on18aC2wUJbChlUU29bpreDxi
feYDm1y6bELFhrwx5Ayyn2UV11eav118HTebwIt2PJ6eP5r5RvdCBovYpzkr6M2KyrXIT40+eEyZ
nsiiVO+KAXWiesaiF/UONjRFwQQEkLA8Fc/spJPoPOGkt9jIHaUBjYo/ndruJ9CXsaKNQJMSWuk4
OlFtfBqJIp6wTRGjyjT8ZArMnPbv7y2PIGorGUFxmnuBGeY88Jm0d+88XtUw4pSnkZ/uBHqMEguE
TLnkA2HZHVhzMB7LY+dKn6y8VJyYt562wk36HKGr5dO3of+vMPTOM7Y9VuH7YigO7zSrJnYoF4rz
Z7Kba/H4EvutZsOY0iQtJ5NNGSqamVI0OHc3KcrRTFRVrms8Ehrwbf6gR2ygUWzreYgYnidyaWvy
8+JTcLkw/J9EaY1dLV+xOHCeclhkk2ljyXnXYw8nFMS30BPyLKy+I/+KW/lK0iOVxIvjFkERh8Vv
c/xnuiuYulN0NgS6RWykSCA+XeAuUrZ7kTsQ4mWMaPTjMY85/OKNugLhqxZ4G57RxP0JZOLw1avp
lS1PHPQWMLyJ1OfsKzkJEUIgc+ihBzDzikaEu2ZeEiKkGSG9tX/zY/gooxD0iNeecD/mRp4jJXR/
ubsSF/DvBXJZvr1NfOorTZAcGYIwdUCqkv+0IwI5klBMt7H4i5lKa4rl3efexz4HLd+U7yXgVbOZ
Vl9oZR/h4TwSkHBWaGbRNykM0DiAsxqQqnl2gVxmJ6+zPARPYRvRoo6hQohMLEAl1syXJHt0pzs3
Daic9ukXVSLCfHMNaS0uhylEqN2xqAWgO/l/fUyGA2OkfL41sgzMUjYyeWU5pE5M28Fo4+CjUZzF
5Ltui9kvR1rTgu89nYXWqUEpxt102sBnjw5E7wlj5nrEXKD0+W3kcEe2NIRN57HJDWfAMYEl9cPY
20G4qL59ixiFH3g8TOVX2FYOVjRzM4WNUldhVlcky58f/E4D1Em80KoNU2g439gQDNVmnV3oLsTG
afJ1XDIAH8/gM/jKizXzUJOR+tn7bs2Wd3/c+Y2H7mC4s3uJTdKM7Lr4ZA8b9ou2Gqsp0QhBmVvv
agJcMTlXPtxDboFj8lcbehtHPi2gullL3I5vdnlPn0U0qAE9A74TJLXA9shXoVYYE3Q66zLO7hFu
A5UKadMmC4Vd+/Cla5Bj/yPO12TE1cJmiQODQ/uQeQkuU6+EnN1Lyz+/3Tdxo5VhY6vJOjhjwrP0
HVRZy8wJPJC6m29o/T8VESBwAzYv046/26HM/W1apHB+oqlZB8ib1lGXrh+hynnGzcOzEb8NDUPD
nnAZQJtICkWHOYm+WfCfeiSx605Wb/9EGCwDWzmRJK64g7Xl7sjQtADY46EcO90LWLCBFSC6PpXg
ArEuJTu708qA1CKjMUSAolBkTZ3dnwmuSrjcPBZ56uTlrwcDNJC9Ov//Mg48Kv2VTMVxxaod7fCO
a19+8FRBAPNoTY7dYtLKCMwY678VSLiy2gtugzrrVHIgo8UFCsEVjWpjaaV6iHbPsnHTaNb9Q2Dj
606fbFmw6koVPABl++k3h41XLjnfrYXrgFuwc+47ZVkFDc6SMBin1RBU9QOvXHQHVHbXn9y4iYxQ
5Q3V+i4WIcBqVdo8nF6TK4YeDkiZbWUi4XsaSEQq0N/zrvAjOk4YKqukoeLa2Bqt54z8P1p/oiOg
dKCXRG4G93BUDS/n+gh3+oueriy/wtXglAzk4qkVbZWARCvpUs/DuDVyUiANP/3FJp910+ppEhnn
zWVw7/idiEGsujW1ECF15hYZ/SalzZ6475f6DfYykgmVnMsoWd2e//PbeT9IgDzL+DYbH/DZq0M1
/KD4TzsknVVim8MrArUBKygWtRiI5akfG2+XfjGTCLqpkzuHWMLzH9teMZxmIAj1tEVENpKlmyjh
KnWQnPX4Wml79XHDZT9YMvVktwRw+A9iookL1qzgS9Kyw9FdK7RIfN17BKw2dpRgma9dgXzZ5dO5
7P9SmpAi7VfCtMoYmpJ5OLEPeoEWZbnvOG1LXywwsZL3mhUnwUH9X7K8Wl0chJadYyzZtsrEX0a1
vW2YFBVjP75KTuG9HMGyVHoSbC2QUe8iphw/QICyIkZrXBr7WX8mvG3KW23bDo99jBl8oK3AIRCD
ViyqsJUe+vyGwfNn3p08Ddoo1mSTBynOvHJwQo8p4ZFBzPb7FFDalwvDzVI5wkO00AIab9ljYwFN
7sm2Vb+9j1C7j0BlT80WLloy0owSsPOZF+4qDgRBAEUBYOSx4NlE2iX8jKA3IvJPnQ0HeKs43Fh9
Q66QiK1wgWmJN8ZVk/7LcSoSKcY3fcJrXiRyx+6Ydm1wKAgJnX34ta58+PT+stZdu7ds3RgZkl0S
tRO2d38O8YX4ZUtxXdVHNXXn0fTUhO5XzpFEmaEqN5hKb8m8gOZxH3gLILkS40HYH953EzcSJOpm
H8OaF/i96a5tEjcSB4RFKHipnjoHJVloRyCzMbLS99txW5MQ8XTzGnPYoFbb+TqYtbhgfpsOcMQ2
nvFVz0a3wt05B3tqYUmhjgHY+WGtwRs9CTPNDg4odMzeGkdQAepIo5LldcCgCVnrZca8ueNOpKVw
Xvc4GZOndNPEqov58FdeIP6vyKdxik8p2LOO5LvL7OkxRcXO6uUamnX+tLkwmeXGqAGTgZWF8VyO
POyWbam3cwkfXkIcaUm+WRaGM4HdPJ5AXeUCf3zYNdyaAOqrmALbHj1nHQv61XRPbkrWX2cRdNGf
rRFW7M+F8bBXVMUWSQCImXFIhZahyo7jui5nzyAFCj+dQVEGk/iuME81JKvw9+m3YalnE19R1atT
2ZbPSJAW1AsYCnn6AGAKYxFs45ZdOQT/lx/vjD7zeFwAKJWy4BI8GbLItpK23XfzXAYnND2Al8wK
7PBstftGusOWgmBNZ+1Qd4QcHpTJdCaBWwT69E5GzwBW9Og1X9etAqnCkRAawvyBXIrupffCKGMk
iC0qMWy1bXlEoOjRlXkWn2kNRMBaK4OXupxM2TUTCNgPyOTO3U83t+gL3NXf5ATIDsGzZOVIjGvN
Fz2I3gidt0AIaXVf/QPUf/Xs3JtYQbEjp1suEjf6+exTmaXH6vPNYiW7eVuk0d7MtID6sbhCY7RM
1lIY5nRhjsTS2NUz7mS3CUbVThzIOATTP06s7WOuoYaHqt2jQI6hYPHQvdDvUfmtPwvBscPq8zfc
IyuavMg/IioAFKUBQoc+O4vwsik5BvjDJCOiCYsp4GlQ67KIKZVxDFTyk7YyUL9HDj3NVgVOJf9j
ovyg1PkURYPlN1h+igkxg97mRk29FPaXJPKrSk8qq7xB7rZY7Q7D7qoBs0Et1nUgI6lmbpduTSNv
DQJ/vdEFCImrxgnm+ZR+zWZfpGT1TjmiRjqFn3vaW16FDAkmEdxLLn2MutieH9+SnvVV9aEsYsWH
eHH2ldB3O+Mni9368vkcA1jXaWM6weYgY+eh38btpuZGPGCu91y3RwyqwVMEctVaq56E4B6XGT75
vqlmzdUvSkC7js1qSdW7BdDQAs9DV5zjIKg4porCZCCslqSfJI8oNv0TtmZoxUyHJPgzWj13Bbie
c8pYbi/DJVQjljLZvfiIlkZhTGdA8+JZ+LgYNmdC2PqlkVsJ0lsH9h1tGdGybSZ2ljxuegB+CpXh
gfLj7jc13U4M4LDx1/PF69rQvRsQ4BVBlMOFufJHHdDeXgXfVhnZkdK3YFmN9hQ5Y99T76zJ+NPA
giNf9EIq72D5XKRPuk0wCZKUT+2tSaDgrybcDljW+PfPMQ7OPTo8YlY3WStL/jq80mDuZZ+IjEdC
u7N1YkPevGo/dJmMAOI0g1AlnBelx8vp/Yx2PxzNLEZ42/il24I6eOv7ndEvf4dj699mNQWs3GVd
iKS3p48qZMC1csNISSDy+wumbO/J0Mya9+Gh6SSSlxhwb8LNNWFYucnUAlXuP+V4cX6ipmZiawrL
K/TXn0ZBCiu037qOG9sCJoWo0+bj95iQjlqzd/E/5WR3uvFEgBPnkZAHFYdbh2T0qhxGyGuBeWJr
LOwtwufdVggeO2F5y/1i68Xe5kNAIALMIK2KLVE8yf4P6VI5UpgD2Uyabb9ZvZB5N9j9BrqxkhDw
lJdipu9sQC4nlwzkrrp9aWwldEzSkWS3660R7OdvcJPwuk5kP9z3y40AYKudgkeIZri6XawFREmK
HBWc9v2g8ss4kFrPFLhP67P6l9vs0Dv7BMimcLtRNpt2VqsCjmLKoF0pTMKeU4yP448X7aGQGJnh
+p08YMXCHXxNINyJPFjKceMrBBlYlp6sxBh+EAYSF4U/ZELsqWORXIuDoid4JSVnwCs9FWtE6UPr
R4xrg4WF6XvCcwlCrUbFqjqe++OoYnsMfdXHo0WrNNgDFaLOZL9fqI2Dh4vME0BJ64FNOZovPFXe
gpXcl4D7JT/r7s6fHgsN/Dptrz23VB3KnHqmxUIgOE0FVptmgmpcNibUm1u301QJEIM41dVdH1Hr
RMTegJ0x3SiG9SCU/OTDQrdfp7K6fIDI4DsfHB3fsoK7Do6STreACeHW4IaPQdP4eL3YpfP/IVZt
f++KSY67BqHOOClWxpcR7sxnA+t6IY9bhaRn0ThZVo/+LYDtzJB9JIzbwMalQKmGQ1qGx0XtO3f9
EryT+ZEjYWPR5lpyht7j1nL9pyLwh9D9yLRhZmqo4yljwboihcl7XBOl17NyMKsiFmFjNkq8PCq1
MU4qffC12mjpgFRpbgiYdCSuDuJglOQ93TUDsowdjW7TWqwL8vEuwTj37GjYjGsnEABV56oYh9Pr
U3/jyTwyNlPYNF5Oyo1hiiKOiAdH02IsS5IesUFaU3/A9YxoIanCsptdu2B+bGIxjSyHTWZqY4d3
9r16N/cyb0BbuzYXqEgIO2pDpRNSZChinX6LCWz5+vNHXztWn8N5qdG6ZVYnF977ZEstpzGogw+O
wn0Y1UGjohDNqlRfu5/ySJVi/oSs/nFOH57PXZ2nb5163hd5T2ggumOX0c/6YUXYU4WB2t4xWm84
MaSBOwRA5i7lNmYoDs4DSUu/BeHghkV6agqdfjgvkUvjVfVu0tIFTCC45UTC6oJq6TFf7oWyf1uM
aQd8KJiUnPvnfn6GaZUxC17ykH49owJdD+65CN4eg+yi9Pp7TZ1PlJboRU07+bN0bUZclMXp2/kp
kUK76Iao1ZaHRiNzMxk2RILKwVNmchQC/nnkbSRX04I6Nven1cFcVIAj+X5/qTGYdylCfSGGCqXF
y5JfK5poU0DZH1JA3x/HYiDigaw+u4wUYIKBBzWC3JFbDWaVshTCsVvFEKfLmaGIE3sgq3mBTfcb
LxiMRXwTReR3F+Vb53f2h/CDEoOJIBPIbcmnglvhqDP8MRKI35iq/z/+rARIkx5TW5B7GuN9vO2e
6nDFu00i2TQLinU3I/Vvt1xXVwceRAq+KiazEAzIE0M6jzbdrY3H8dJ3cza+jMgULaEMpOBaoFVP
ABGjAhB5QF6AHe064X4b9sLzJ7e+9mxqm3bHU8pCNDX0YOn3nelacuIEeLZKsdsrSZunfPDmmb7h
LuIZTxJk1gj8x9xjw1OhZ4XIanvsy/vObbkoM4b43HcAubRGxcYtM9wVXtm+pkBXqkEBJCu7Bd6y
sfp09zducdng2vJAGu4pp/OIEHtDCwTGyqBYje3lko4TLXkZk0d376HXWrtWKiEmidXN6JeI5HcW
3hC6Fq6PsaoaB57F1cn/CfArJH/T1z1gIlfJ/s8nQ7uePq3pmOsfBtp0PWSlAR04PbR4ewxA/T5R
kJhT4nf+WiXojCitwM+mUykbChXcyXhkz2Zw+IAIVpLBBAHQ/Ov/Rbtw1Bq9fmv4ZNRI6LJWx4dD
9aAGBOibOpdvWnJ1J8XAYOC6u55mtgcVWnsK782n084DA6I120gSTt4kenTR9WbgEERtDxDW9bRi
+0ZgmAt28pRAiyO6LaG/J1sl2n/2Xjc4FrXsacX8XSlqJu5qgnINqDR+C1QNBwGApxxYS0Onf4E7
YY5+Frj7FCnoHrjjj4opOEI8EmNTFut1vg9dFd+675hjnb8vZ0vk1lYgfwbUu8bGbwKKLha3Jff/
LhUPlQi2562/4l2vFepGYSPA1kozu9PAaxwBSnl9/afrRLtKzX4qz2wRo5B3idb1ELQ2b2D2hoHS
LnuAQ0p2DKfrhbSe1mGM77OwNIr+8DTTfGBMdOrV0wqe7/8+qNJg1w2uebjisN/5TFbqjSWgTQGQ
nBiWAkKMQ2iIbrZzvURU8YZmfAU1jPv9pHpwodBruEvFjlTD8jeTQAgvsJk2fCpMHktcT+/HX10g
x9e76udmzMzSN0Od4cJfkzPg9lae88o94/XaBCxy0l4u7z5tjTMQ2vwDNyamjgixEPdT6pI1l/6n
RAKUFf+H0kITxGHpo8vFwDp1lAAjEIP6BUX+eQbhc95+6hh6nLaSIMwzA8g+rRXdeqCyEftghkLv
+bxAVFirlG4XEj1YPNyqYbLUWEJK1HfGbjNiyGD9x/Hf4p+5nep0/NljiIUK4sBP7CCtHajDmshI
bi+1Gx5cQXFym1ose9EFT1dATuztV8u0DbXihy83VLeAxX/pLky/qiJWlVYy9IPPy7gtJrkfycun
vcu7Peel5ZOKEgyFCK1khgmBM72Fbzxzwnl1EpcbBhQSKLf/N26Gvm06T4tMYZNFFazHA35xqsgz
aSycZERERTCOBla91RYqDbYLLqCVBBt0Z7XoiYPNQjartVRQE7+Vtpq/IzD6xX3W9pUQmJdE9aIN
/tim5ZTx+fox9hhlaeRJRtEIRbfViWJI2+ylV0qLSZx1mxz5zkEPTDEIwOQPeNSpysj68ScHoWY9
5NW47Egx5QV7JnYYjy4/32iYqctds7MiBkVttESmt6IeJnN864PcXhUkl/UlyIGODLnrDF3mgzPd
SqyEFSA9ZbDudC84RdMzVA2edRi9AFRr2f5IoTvrqFQVA4YRQqbWBbf+r/buuACYkYVSzEebQ3SV
xEwtAPddG12KeZKKqCw111pz32CEcDE88GXc2DaeUx9DVnUe6IC27RALFJNCE+Cky94+2FBFSRow
zPRtTJTyV2C/7U+YCqI5ZUM1oJBjqP9TUjSlREFEE6BSbsRFKRNA1T7+siwi634lHewe2+rofA1a
cB5h131vbpH+EVGe99oRGw0FVlaFpqzAgEfip/LW3giZfcb1Y5g6f61t/aIDWRq9RdI61mrMJNQW
p5j4a+IOgfEj787YaN+/u4VcQixhYDLoujMrIo8RdOKFBssMeFA4bxh+cXSRiygnTRbZGVKkFN7+
v/53uLy4EuC+h7+rTQ0d1wgtXEaueiYeG5eZEKk+KCRzBF2u1mtGKgDyZveRlYYH14mWakJFVAu3
AQWuo2G8vzq30eUGHZFz5IV3bKJah07Or0iB1Mul1laeQFiYIYKR74XG+Fn3lgxq6v9bNFvCIJCG
cBuREF8cR/yHwrRy1SkzNNKWjhx6+7nR9w5nTHZ/lFutlaQEYkFqEqu0nu+2boPpLLrGuWE74sQa
++X7Ri3FlwnatAbj0WxbBNx65J7BVQK1rcManwXXNo5z84izrN1a44SrJT56h3Mm8HTggg+dlV76
pBwuCxyLP5/j+36hxlZc55Dwq/dhmdPG8AiU54NICkUJn7jG6E0dNFA1lIYHlRgSRimKqIO2d7s0
1I+0MPN/flinU/wKP60gh8mbP7fN+1htGpnvFnTi5B1S6kH8r9890bJXXve/XkHig1qUz0XNf3So
dG8IoHAMHJc77J0eLlLVUFPbF+4dEtkr/7+1EbqUP0Y4kn4TzxO1qDMcDTqooc8rOATex8dz292T
h0hyE2sxFwE8zsWMBgzWMBEa5/OGIOfKXVWoiYnO6LsnR2pgXZdr5YOCyd2awymLsps0HzG76LHo
N99MwBwQJAOzDdXrFux8+3f0tS0nxib12y3p22+Ezn1P1u616rMv6XpHFpWrN7RWlryjH1KT1tqT
c+QWDFfDxSfjKQp7jSinXLDeotDnrIfgc+VlpTl9xJjuTk/ttCGcviPZurdRg3D2b0lHSrCguRt5
UXfRiqCnWgklN/e9/FWlBwqmknqGLTFiKR9xPTF59PSG/NQdi4F+kKzwJWDR/LRjiWmxQZfFuB6L
r9payfKAzJ4645QjgUTfchasw53z9EYpGUa6r4Z/i6cq2tyTDkkB1EQCaVLHIRjcBK7cXq3fGQDr
d3hg+HTI6JfhnXVivCRhd3kYo92HTntpoZ2x7Sv/wd3BlQ6rF/CK5e2dMB0O9gfZQI/S3A0guFiJ
6dtmAXG4ZQlrCtL8Zt//x/xTw85EYBfB1sox5FKTNPP6KGSmXVVpmP8dWmcwqqeesKCdkVk5XveO
3hLQiZ1NSppe9Vfd7O1SsmxyEPI36/F7YrXXG1377/0YzJAI3q+TylP55MgA/hMvWF/fCwgyyXGq
fkQ/Ky9Atf7K0cB9GmiYq/+HYMyEnEHGUaS1gv1BHNltoPpDqXIQh2Q27dC3aydBQLpLYG4147/8
SmufTQpFBMD1Rk4x8p3qd/i/qQDP4RRR+IvyKNM8uAKsjfxu8IeJiAjdf0wWfHj5YL6xSLc43Yvj
c//zSZYJMIihdPgMQjO24plUQQCOz0f9WhGyCh8btyr+nx7PdS1XdwYdk7fiMQJAIvhVV0KBrjJm
pWKadvdIqWErWN64hpA/tDVWC7b0D51ikOe0ArgoClwz35p5uW/0NiP8/J8qo7KEBspz0tyykX7E
j+GqUOvBaxYPIKqfg/HMMbvYiSTWa7D0keeEqatEngYmBIrMJKlkwFjh7FnPNmoaJwJTBncjh+Ql
SdSwkQtL5QdbhHxjKrGm0xu0nB3XOuZ1yXsfVuw5k1UTOfNa4v2HJhMhWxOn850IMycRWU20T8rg
+TUdpsDQr3EEgXyxcAcRrdBEGJm7qjA1JcZn/d3UK0yyYk53I8/HL+OLyUVvxGzI7ORQ0nwBNtu1
28ZBRtgUx9oHsQvAnC+2QR07kC3cnqZ8PXxRpLj8JTXVBA10SMLnm33fjx1bjlm50df72YKSYD2Y
wfyPqnEcAy8/SxqIesOMxn/P9P7d9aMfw2WUz7n4rmoLUn6jA2sqPUTnqMyqFINWixHD1MWWHrq5
mYfqj71/mqWA/gYLf2n/wqQq6NmCEysf76wHKTKDPeNb+LATDAWu2xFB4zTt8xaUth8mMfWf/Krn
BZAcNqlPYtGVDfv3Q/eYCZEu3kWvWlvIifc/S5SnesPhbr3S/NKAyvHEeJHJCqJmI/0AP04NQpen
4frCkA7wew2FO+PESiMzQOEAEKdzxHIzAeGJFwvBPxl7j9t2e0vjDt8Il8zLmO2r9sz5OtGp9u+U
AZq5IAosZ2cEIBOD+OUO/J0cx1w1iDily3YBDyCsgH5+GD1ipClwDNLVCguxmsccP9hBPlVgUjHj
hHgoZDgKqQEAhZgL/d4MxxoK71Uo15A9Xk7+pzSFWtsOJHaOnbbEXYVa0yo8+iFTlreMsdc/Grs9
Etyo0gmkMkwDH7Iu/HR/E6nH17Qo4fg9wCQpJj+VjLQYffYXpg3SA0/bN6vdE6+nsfVejClsl2oo
c13hwofmo8Iq2EpxvJbBVC4HHyT6Nja0g4NOsOjfsBV7nj9FB6qNeHAYLNcmdynPCdXMq4K98jMA
HfVV/QI2tQRW2vRTa/IcU5I4Ev6YyrQZFNGNFTGLYjH2bd7a7QKu7rKI683ScADXet7HT1jCQ/Vq
P9dfAn+l8CWIscWR2Aj4R1SjLys0wGwaCFdEtEwa4qX4UZZEU0WSljjPqUAXZ8jMNDePQ6CoZKUF
4uSuAmo8Yn7Ew57gJRSe29b/Z9rv++2CjPhns+cZhzIHmGxxYSOGyllnj30DWR+Q31JYPImqofiK
lu7LijnMH3JzWOC2jsCiDGd4luvuswseWxrhFnPQdxrXSYEvcw7ZZwYmCi5w30ioPrLmBdgCzQgq
G9c8Q1C3g6O24/bCvCf9ZHu4HpwO9goKummqLi83IG4PZQ9GI57zIJAd8ywOtamJQaKqp2IYyp7y
4nl77UCNmlfA5X+3Sj0F4w2QjU5k2s7NYb9o6A6Da0Kf0QzKAokwsbPs89T1Cp7YeWAeZJ5d5lR6
wXsvS2pp5ojgFXZLtO95QlyWEGZu/K5MYqdM2vrIucbog8K4+qC35zgVaCQGjxPP0pMbL+aLOAzF
zEDlpqU1Emt7eFlWxXgIgwlnNasDL0/Ih6E+MH91oV+D+QewEEN0+xkmU01FA/AIizokSyuNEdf9
NSc8oXbXE+5v6CDTzQ1VYVrEXHSsrFS40ppj0LkDRORbgJfP1ZmGdbcRGvibQbwRL70R8vAgzvdm
NT0MX+5knxrAt34SkPg9tqER9UkTo+iK7bGKM2Tzz/LRceFO1+mMQ9bJztxNmkjSNcB+1iXn47/x
B133DGKE16xHVRoZrI71eE+Bh/EJ4Ow1xY7Rd26GfajxNmKFrp0RNkZD9yB/oUOxQzJ8bkxbuia+
6zMI5blkC6iBZ94e0wZXNme69ocpwX0nLAbuJ2TF7zB9GhdPeFIpanFdfDhG7IXXCFvYT+wjBwJm
r7e5i58hFamecVlroFObx7eCgA39+BqaEb71XZ5KpgdIuevCKfoI7yBMFGO14h3gPSZ01eoNDRTs
OcTZHYb/8wIt8qSoUes9cOv8j28gPVS+D1XzZNF3sXsrg2/nof3VrsKSX4UEroYnQtooUDH5AN1f
KqHcfetFnCsEYIqC6kBNIovL/+PKEPDAKV2BvwEezA0viEVlyMkaLHYVtpmCBeiKk/H2IwUNhAfg
WDAgCY2p2iiOM1PLCEOw7XBVk7MjWk0x52itRLEbnklkCE8ytn0N4w9Q+NL2SrikZ3CHcwhuwWAh
XDDQDUCL3cZm9OXFMUMJkMpg0heHejd9Wkuc0+A0CUW3YMgdBLttuSyEoyiMmtc829u1YAy4iIuH
RK/ZOeNIuFM7iaAfa4BSoD3Bcp42Ejm3oG2OO3ybRd4HggaG5d24esWXpBrdxiXy/ckI0C2GJebI
P0xOt4E4BDXfBDbL0vs5GFSvGB7PYHsi1xfvndUwiLk5Qb8ZDia70jFcRPqvYlsgHOciRQGiV3Gw
YWZs6nG6W0fN9wguAL4qMrmj8nF+4tCVSMXxKuwCoSVfYG+3VQV84PYS4unatQHcRKxT9Vb/m9qZ
/xt0wPZgt9zctC9mwCE5iEDh/YtKgwJYWAR+ZpCSqP43DbjPQCgvOIVr0R2w3Wx0Wl0HvrcA+YK9
ttZ7PzjgSA0N26p01jTV+ac9zQWR/OoHJpaZcjYzEAIG+Uqq2K1iZ1YOVoceyeM8PHoUtlEbru4b
6s8HbrK63qHgQlSu1pOv0EKKkyfYKXX54VPXo/+m5VNGOA/jczIcq+jRnuskO1kfqNKJsnGIP15w
HmWX+lCfFcc9dr/uaeGL9tqd+h48mtmm0I5/BdsfbkWposAe63VEQZh2G/Gj6K3T9adfKXbr8RmG
vBwp/Wi8BUsAD/9UwtiyM0NSZ7G6m3wT3oRxx5A+9eBPZjcDo8fOsRK2d1+juoO1MUdu9tLOghmY
TaFxJSeNV7YljrxjyUBUkvTvfwz+9NVtyx1WFlO67Ueq1A3JeF8kNVwJFa1y0Dt2A01e/1WeSKyd
m/0BCkG2jy7TK4mNTPBfc4TqfrxpB/VfgglAwiLPWw2ZpwLOGWKOQbvmMMRgSpsGnb4GDwiUFrr+
J7GJaApvV+46Qxzd8iWdMUKM3qE8U2iB7PzNyB8gJw8oQMRdSf74HeJfKiqGrFuV0YPu8ij7pudj
tlfurHXDysLEGkHYObrqYCChp0G4C7scoDcbnOnEklpOwg9e6LxcWmA0tRTUNzJHUiIe2EgfuqI1
qsM685i233Uqs1SercYUc8yZVmCSStSZ7I5tMOnm8X3snKcTk8xZinuRNL86XnUILIzBAWK38eDN
uCJcAnb4ETgEG+ykJlL3PiJ9Uj6nOafp8NGN9pmg/tU5k8yh5SroZe8wDYGV5UBujiCEh1rDQKjW
NURziwOvxnvH00EXDi4QgUDI5HHgMxdepxn1A3mtmSbPOf69TViGxUZ30nFjSangQVaD721LsFuZ
evdmYgqPZK/w/2C5rc2hM7rHb8LXiTVpVFpHkqxfnNizU6at5Mw8Ui6h6wIyXReGzUEAFPJ9bQtq
oLHq64KePtepB9+Mp5YvQmBU6+p23DD91xyjR7GP2hb09MEoC1CagluBj1NizGXVoFFWb2izCe3G
jJqhmO3aasNjBLshuNN5n9zdNsFSmpAaTe1KWU41Gcq71Xsv5dyJBU0O+H7i+UazpyQdCULfnc2d
3IspYV92A2FE0AseY2of9xc0yhEBMgcXBmXo1oUulRvDhEJO+u906JMBtE28ZdWM/Eq2ZnLYECkV
DYEhJdVeqW8Cl44WN8WW1G94NXtrP2RlCVQw76c86a/aOkOZgEnpP0T3wfW9NJL68dryrTzrju8L
Yp7ZGl0hz5c6yXgsI++Xb5y0WVVwsSLtt3gC6iyGFmEwzA5I/q44qpnn00ghwFWDotnKXsdJ91YW
5mkevfuJc5JKYdFckpUzxYoGlOxW2O82DZ2Qx3zTZYeu40x5vqq1FmlNriBmXlcpD6VvRiuSUBqn
a/j0duq7zjarSI4WqZJX8pBVe6J5Dxtaln5dRURfAEJnCeNKRz4w3Ub4q6BoRgGDYP+GZboyJMvb
XH/JvCjCWyCNiqGO2bwP13gfSjK2vW50d1yCidVCH+VYDOj0ghJvD3wojkjBngNLs96p4HfEo8wJ
y5nSPs1YT3q+ZyP0CoJsEcUY/p4yjjbkj2JDp8qLQRwUK6LrUqLJIARzQU+lP95K/Teo4GM4jhSW
TVvOELu5FmrsJOu+MqGJeTmzHxIE0ku0p5DKS/uAhCOAo/dpgZF9Bj3gybEkytxBUuSfSOZd4mhR
c7E02Vp2IxJ3kY3lMJqU4lRa6PJQImEs1A7ywMu3m2hfXQNTfOKVidBO1OQwLcyPhraUnuW3ZKmI
7BLlehhQStqrRGCU7b+CGYtxS9aRjODobOJPuVwjpYxcFp8htTXi8T3GrK9mO1sohSbeshVB5hr7
+nrfst30IuGEI7Upjvk6nBHgSAL/XACGEvHsoep6fGrvP8utLfhNvq4Fy0Tpc7ifrtPqFXIaWjuM
+efsfvdWXD/w1K6LxCrgjUswF8yqeEwZwe6fLKde9z6UWAH6aKJj6P8tXHIk0aRuc6BIp7ytXG0K
4NjNgPmW1OstpjEQvrlhdwc1KJ5+pSz8Bkev8qTHu/OBwlCgeBQwNjuOTOsfhEIJ/5Ww1LzObFM5
55+me5I4LCMiM6+GeIcdO5No5NCZyzzp67YhOv9l4WfBiuY8Cs7qg20xTcqFUF6YzdFv3NyVo1c1
SrbJrTAHaT1OeirIaw8N7703+2PabJczYfZ+87J7F+0qCv5HAjFNx9p4DoN966bdFCNH0BlSfhfW
PjfwkLIqBwWOPbHBYuI0ZmjxAousieS8Mjeuv2OhWuVhRpPJXM01N0hCGybuvtnXgYXbnroK4A28
a4YwoZUukQOwOHu8oUa1YwB71ipBWJ6tQGd8M8VFKZs8rcCIGWZscyyGUJyRn6BiwsQLTW1hzuBS
o2aCQNdbTxNOYKtPnZI9LTam2nrfP+8U8FLw76idZHU8/El4VyO2hhGJ5TvbopSB2LOFGMmsmKuN
YVVbygYmgvOmxhEWnXe3Vb+TAQWNo4m62aOJKH0TCE9vXsfTZnnlT93Uo8WMbBEt0KCshCCyLf3f
s7WiIbmHD4Hnk7mHFVYBeT+ZGcY00mA83rYbTjJsNuK4vM+cmVs0Qk+jIJ20C95pNQZLZSGFmWVE
EhFhG/yVvVCYdtn5FIirwELiBoDAAbt19Xr4PbWtiVNhgqbqXdA2Jzrxdj6X68Gpp+IGKdKbmZJj
P+I2XgIRq+qS2fgd1f/rXvz6EEaCJUYrmmsPRmgriA0McgsIUQQdpBkuAVcyTWpDyXoeNTZ0aTOZ
uF5XY1+AMCj6ANlLKbz0hkQAh/ve5PXDAhv2B/KweaG+uSahHDf0NtDMV7gZCx0loWX/PxyOfNMm
uw37J+9ejl+UeZUA8w3rrVVeq840NbBNBTix1Qo9Gx1lFcyRM8RJO1X6P7cCGWp1I4U00GF2KHVx
3rldKL5yX204KxentT6gTWxTYaIQfT20gE2s8yBA1b2931C4lvKB1AYAbnIrldhrmVr+1Vgkz9NH
gX3FjHTuJxmF3h1EbTAUf1vM8dzjDd7PT/wUFa/GfdVxAtgeZoXOKudy5ySVUF8ZXstQdVLwTZaF
K66owy+PjTTFQTrrnShsjCyrjqgzd805mE65pUqn0OFv5VIu9nIWuPYJJ93ib7VRtRBQipNLNRCE
+VJuoftv8au9160oSBsHDX9uXQAMQFoMTlAOfR1HSVpXfbWHV+yDJH95k3srT+uZx/lsCUjj7fad
K+j8Hfx2XBHjXZQw4hdMUKJeW1K59vIgkcs+lztyPfbL7hfzTR7CRJleSUdWKG3KKP8ExEiMxZLw
Im1T4FUGU9q9BmvlhNYUb4bqiYZa76ZpTYLjUtGgZOz+Lh2nYxWdh6YWiJqiKt6n6TdI67+VbG7W
GwxSwIMLdRmHWT5o5gBqrCoqxkAkOAAnbczpKMZKle+u6cN5dFs8hOpHzWHQIoEcWw00Kn7Mbpnq
s18gUbVBJQeef2mkoKqvDNnBwjkaHmHyrP7iUto2MxlA/DrQc77jhbRkbE4MZA2ZzCdKc9C/rWfZ
aVN2ismHOw1L1xrZerTdasKzNr9r5v5zI4ROkxwExqDcxTRRXzoBWEUuB4Im+tQ2buWXdbkuBuN3
uALAmVF+MaoxOShsrjAYmRsD+SbXCyyex4YRCT41gM2T5fkDCccR75o6xZaCs7dn8Yhmg5CD/abl
pi572jfMGp+OMwEifL3BpkxsV3s/XktLDo0/laphX9ud0l/iXenL5XER22FEbZD6m9DpkSUoVeRO
HOj842J8XW2rFdmcQfu98ruppSkE3NLOd9pQj0ANvuz+czBMkFzkcNdtl8Isvz9LFByMrBHKiV2Q
9S3Qj2/XCFz3gXzI22PW2zva7etQJzOnXLisRLDiBMWDr0KG0pF9ID39cKKfw8Hky1dQ90m/7Qsv
5JmiDO4n3F3jAE3UfwBCGaQgM9F6CyKMd7ZePT1YfaruwPTXCdeOZWT0doVBgIoApTlhDhBHtyvx
1jEJIs1m62Wnbu6Hl/w0x0udwHxrhglANRX4MNbjyaZFacXKWT8MesuFmYOv3BQO5qb39p/NOMJh
XYmLKeV6YAaaf1R8dzjYi16Avi8EBHmP2yqgkQmP9ivWBXt2d18UVUtZI4khGUGov3asLhGMVZTT
Sycp0/Ec7Du50BIDK80pX72v66YYMOog24icx7KZSAkM8cb/OzFoA6Uw0BibWjhxMY+q8cbFsbvO
TUGNE10e4sTmSSiaqPBf3VbC7IdCbnamd94+i2IO4xnNlLIb06o/lWcWGz2pfzV6DsuE1GQ8dNKz
JECxe+ior3/k/ZG6nU8IaeuUZ+hlwCijNyRatnRdWnIr72IfEcXRXwsFAQncjeOyAfVmlYTtoGhr
OphQEQR4d8RY95lANkKMhLqeU8JXMaErSATeNClvP95R2WVR5TFzRNaK3Qg+iV+yxRRAcjObZfM6
epOVzUAhvMKSjJjcO/48gTj9LFhv8jAhv63c7FAJNcVrlAEcVDAgw6HaVyIs05bGfJRNF2a5kyBS
DqAa91pIHNAGRMVFbZ9CyiZJTfsflLdE8yK5ZddvthvtP5d/awkOeRV4mhoD2e6QPxsjTl/TBVhM
aDGtKhbd5az+dwXtvmMN/U2z+HKMlmDjJk3vsFENVDzIVO/hf4X+XTKhvRjq0RWstB3O//N4FYkY
wfVLpDiSanYOtlEFLoEm4IqP05sRmMxC5s8mXfwq78ki+f5SzJIlykho0zS7nA9XXtHZQ5iNrrS+
uRWlAMShPZInTOrqPiZZ7hpqK7LzfPXvaaXsii7tE+HNFdjJuyDttz8LSTriBxYehhEMZMYRsgpd
Cj5C+yJ06xVqmxZJrsH3jwbPkilkxo2YMUJZZEeXzKkZSS+CNTAbbuoZdmvL4d0xCKqQSGBIYfO+
FiiUYv7FmTdyZZMPpZWoVFRtv5AlDk3SF//jW7wRPbWIUokQ84/Pytp6aIU9src4RuHT0K8Upqs4
iEsdgLEVoLicVpG2jQvSuxjW1RXh5xF9rA4rGLQaVgWzytjnUlJqD3SnLbZI/YF6HQZC2SivWxcF
Msm46FoxP04bIT53FhZ7kEvkox4lNtXXPTX2iKeI9oOj8HC9D83gQtWgBoxymRRQG8vD8i2gZJoL
UTG+QzWr572Ieb/CiRqCo6ZIGDuNASaK1Utca9C2AMYlzHQHqHgOyAMJUF/nVCOy0CDq4uTJWebb
Ka8A1R4WObN/qqF6oC9V4c1PYb37XkcSo3X+tfxd3f+vK6/2tFvdzaq5Thl7Uw6ZRTMEYJyM8D7D
aKhuaAqB4CPyxI/qT+VC6YdHAGDAOEWS/aqNcFJGF7jbMsX9UGOrc7157jD/8oKuIiibCIRiqTjX
mMQ5gttUtYh15zlVSzACvj1ZXSR3ww8jJ3auc2GfqG9COVWrqkDqaEHr3+fMx1POucmOPAySBMRb
Ux/0oAUtDk9SUpzO3IBFby8OFLLJS7Zd0X2rJXVh2z2CrPOhaqbDT8nwN19rLwnjkuH+PYBl2Jyo
h53N3vnFICY5WxL/bNXnKld7x4XBU6Qj51LOmoUhf4oaiSCQBGnciw49UQxmaWcJHpXubQTqofmK
hV9ZPLfG/ckrXxXi+WdeKsWWDoyBL1MWlfiRHvSmqpjtQO0NpEYebnJj95qU4cwnGwVaPyhow78x
biYf3iojS4r7jjSraVTJYzB0DCwIyxKqLk5MFnczNXQxIXS5Fy0qASsdhzJsxzRzyLUyPXe6ENy4
g/8kk1fgMihFFcw3VJ3sChlRd9wffQHgB1UcTj2ERMMp3c6lMr25rP+nKxuS/dYaBhyU2ufRVI+m
+ZHDlWlq7X/Smz4/OFbFE2GviUnEvpeP5zASKRcyrEq3YfEc5j/AZjfORgR4VwRx/mq1ma108DI+
sHMS08E9KYfbo9EsYJGw5+ysaPW2UOOS49gnWb12Is8uF6ewNfI70XQAMGH4Fgn2P2zZ5EovoACA
aRWC1Qcx+Bi6gAHuTXCaOUu9uSjmi0w1YSIC0EKe1sFwACikZKtP8DdykGN7r1OpgYjqiGpaGrW7
FjqI3YEfgVldKhjDHrQ2yU1l2XSnnuQF92jbaNPevzUL/abnf9Q/35pH83uZQg/CxLliPpBTA70g
L06KS0IgXIeipxmO7F+SArW4iN7SLvYk8tA0OtNTv0cFLYzX3bSwJcakBTa4jhC/OFv0SWwUiF3b
s+LXAM0izX1VYh96HyApQEl5hYB2xG9H31uQ0eYkli7zSy1VlNM6/5rXJrV8YVI7uFkLk8wjDrdS
gfB0wthEmXD/tAAgck6rMwEn+nHI7zz2plB/EYkoXqW2MsQRHNmrZHziZfsO3rOCTDdBJ+sFAe3r
hU7Hc30pPsbfJfWsT48miCG6P0BE2Qj0hznBSzCevG2MOLTX130T5zsCvUmxxQKAVhiIecAqNH/N
k7nq94+1D/kWWiSt+GdExKgaVYlSQHsIOF/jCAXgimulEyFdP3BUCZYGIKzAfpaWTMpqF5RS06KJ
36v0BqZeZW/xaCxS4klyQdzIKCix3Z/knVf+4vw1Ws2odwh1Dm5SiZzNUT5eh84BZot6blT6KA6Z
iWEgycQ/MSWkRFhwLGuMBMefbPXWa25BR0ynuODynT1wlJkCHj3VAVJ5yXNSvTnragdMlV7EIiuu
uB5UMDHTFv5ycls0rIdGqy83iSWFcyCTcy7NRtgUyf6WbSIgQQ98Td4K8le0DIZi551xI4ArwQ2k
/WLsPfTkrS2YrWMCXtkujj7OV6RJLJqXEpa6dgLUUK24CtOlchK21zlWaQrVqNvBHzsvpgJd5NA4
waHMYv6C8/jYk1eF+cvWsLoIX9EzmSqJ0mjYTOQF+xl3DcwoXUg7ReKLroF+HuVquznFTdwpDHnu
TZEPYHS7bmQZGGwBBBJHBIn9/kJK5geUdW634tzwrGmSFG6TgGzJwEodnO9laOVinZaflTE4pv1y
SVLjdrsjfydwpZvKG6iMq9g6cMhZyT4wT5mfkuEzb2rHMAyb0sKZrySsz0TUC462s4osaCsAVUTK
KrbLR9x6lftGHGv4bslKC9hGCP8dfJzl9eNO9xY80Oli0gjIONX0g5I2FQVTDHf0mU1TNR1AmpTt
Ms8cjO5O59rVpoJv92zfEGI87gXCh3+mmzUYYHQ2vfbS0soKfYXru8QiRD2Bw9/4RCUeingwYqHg
dN27TOq2YrS95Ifo+jFdpzwG8GrxopGkTohrEhFYFnXyf2dezaBGh9bgDToqGhKAGlw50ymoZssf
eQ3b1d/GfnvleUrM408OcWb/NWoKTRJfRqOo/URUb9xs8lf+nxkruGslIhqAnO25rcsBIXgaGErt
X4pCWfM5S/WvvOfQer9Ig3rhlx4wSuNUN6uJtPF6xdZBt++4muITOQuDEaqVGMvwNwQvmKuhEv7I
GPzzoxxY5OKbdxxl8SVPWQOCk4UYjTnRjBE+5+55R3jitFVhY46efUA0w/H7QtiApczK6J2cohIp
Cd1hLJvLCNSKz5V/9msnnqtixJI771zVTBwukMWQ0tpnq3EdYJwoQthrhicIqdgLSaNVAJL+L/Ku
kwPjMHm5d0iq9bmokdr8ce9pUujW3Pae6YScHJV4PRys06wqKrNRRqOWg2sFtrDymuicbxJA+s4f
E9sEb4/F3B/VomejX82sB8fvjICdBXw1tO3MjBhQ1x2xboMdxNaHrzph29UENAqGf/eaoy6+kURO
Hq1s4k2lFkLAEwwWkXmheLa5SFj5VAJ5wCIi6+DzZWq1N01paHLzmBmHhjJqBAVL4uKSmesIRNvj
b1JDiazSaC1lOYR1JXWAX+AU1Rz9wujr6zcU/cjih4kQ1Z8kJc5zHI3k1IyFm8vz74NLMgPgJe13
/4pWiVdljpiFm3Mu8rcEgLwg711NUXegJbYkS9WjYHeUNpLJ8X8eAV2g9NjoQ8SEWaW+7FXfO9vI
RgZfpqZCgvMTMGqbmsYVcBFlFXgnrB8wnkQT7QpJZ1C5lvvn2EGxrg0atrpwl5/V9IXSUjnG1mOz
M89pGhgQb9ZP4VT1VF6E9DPImZNkzAGMzPDPBiKb1vorSmzP3q4XEkiI5vm3qdQ8ROpO/fWNr/XK
gURUf6FoOo/RQaX81eVBatQWzbL5XPXRR9K3mMIqq8sXBc3wdaAIQmrtR+I22Y4uTxDmWpwirORa
4IduOxHWdHsEwGWTocGEZVzRqYKJdKTGcuz/eaKJf3UVQglOUISDWZf4ZbzABYttoGPkzAArKEKq
hcHJnL/LTknDZo480lgXsPKN5568rvcHjnkDa0S8qEIMOVZNdNRPwn7hmR9NgOltocgEU4yc94BN
KF7b5iSWp0WvJbJPgEElbwyu001xzEX6ja2jgAXMW2kLOe3Y+p3t1B2ZGQG4rXAk9SI8q7FnNdXn
zrOJVZMEokRPO9LDQnUKAaOQBjg1yztXFAwKynr6y5o205Omp04yiLEOVNRFqZQ/gnbM6QA0MjRs
W/FkE0HNnUMJY41IEi3ogRoua8oBBArN3p2dtRU9aL2Pi9FoTBFNOlJdCrU1MsIbNPaLQZrIbE9Z
F/mqm704s/ejMSaVo4v8xAdFtlQd5yAu+tjfVmAhl3ygA3smN2VLLwMhsHtPkDCupnEOrl/zeBAA
KfSFuc5PM5Igdwj/SER1ampfJqQFoqVKSwbf7478f/5mmzlqzICo5XtQawwrSausuUS+8yW8rWa8
eAuZluUCi74GOx9OtRIROLgllUxkNLpUcR3eH3GD7LlQepYoEkqHm2TpiwpvwjBlZdeXAzOq5ial
c5hI0mCwtsoQMTUylRC+8YZ48aBJi+4u8GqaVO7eeSJdsQPJGuK0TUjfUCZE747NADzNCmmVV10R
2BwviylFvyJ7p75J8P/jteSErhEPep91ejnMKSUgcamXR1xyEY+BjPXnhAffclyjmYfo626ugPF2
9rqro7I4Dwarmk9UZtP+6eKiewT+jF57x+7UyoqD5aO7zYB1qRHubdssbzC/7+uBqcvyE/sa62fr
1aWtVh837bUV3i1JGPb7bjUC08Yism2WDCVhChl0RNiEVOvXi5y1nX/dg+DzQbrLDkpLyxCcvz5r
Vq1h/fXQbMIlYIthSWuUFKoj2J75jvyE0DsoUjoiz1aI2Rn6TeoEWpZ6gf7g8C+svjyWkFgx8tjE
6AZkRjiLAgmKiQwINmJCvMWKes/PJETmI4sKaGlBUjGn8cZoFhVCecQI7x9n6hIPkIXb0E9Qppk4
eNTr0JbhipwpH9Sbf2SbxNNk3hqwAZs4Kf9DBTM/JPNoUrQ1br3TaSvhSPVCSvWVgyzOnYXR79t0
QIcg6IWkEi5coBrhTOyqUc9ij3tDpGXZWgCZoo75N3SYiUq09VKRk+OvhLWNTdgIeVLBRy+uuR5x
yueaoFkiJTmRleVPT705EYvA/x7zQm8sVrAjbLlrOGd1EIqXJ8GdI+A7+EgdS692cxrghklWhYgy
MKyZtBj2Cj1Yd9bbwMMlG6wI40BisJxv4eADEnYmPveFa1tOTMHgPH5CMzYRc28efuNrPLzVflTZ
EZ9bsV3gROXM/fs3/pMg8NKtfXt/svPY05obGfMdBev3NF4sM8OGpm3KvyIHPi1iSJD68oX2QOyC
Js5v1ND19BKPTwY++CREpldi9lY0+hG+RKwtElmfFkdzkUGkG2QWJ28aKgF3l901J+vMU4TD+QOc
lGHBszJ0tEZ6hxQZ8cb1jFk4AB+IoEYXw60Msc+4EQJAy5No6Rp8Uc53OuidxZ6D7G1QVKSuAYWs
6/B/sWQ/QN8PtSBbjWS/xx8oa0L6p//Gmn0fRknv0VieQf+UfI4apLgrX+RLVychtoto95oi2cyc
ytwRl2BxjhQAiNTz7iOrD+9+DwohAe4ACoj9Up0aHvX/9gMpQ3udqExbkfdfcI9cqpAZi8vjLeto
XK9Lott+PK/8YYD4qHzrfs06Slbs7HydeTG6ZIwQzGLenyYT7lzcVGfcu/S/m9OrAvUlZb9TMq5g
faHSYMjwYbH66VbHtueXYPOTQgPH07diU5XJED19GhBRhG74gIg1dFHmjOzFetcjuCZSvBQhuIhX
ULpjxwbzJMyILjWUbBDjcobVptB1561fKhRx5QdGWUe+sawDRNyfn9/6+ShKBOEPzs8Cjc6QFgmA
l7JYZHJStaqIy6RHwZcZEJ4DW9XYOmdnTCN4qP2hBZfb6ulMADDVOuFQ29GZ5y3YVcY8lGOPLdwm
DW8tCT/RkV+Zf/124ArP6UnShGKEwhNn/FwNrer9qmF+EMlf8aWalNVK7Hgg/gHUQ7Kq1wp8wg01
cMwDqNz7L64ZPK6rQ2W/cfnXYvl8PRMj+hsVNJEQdUbT5pRheFr/CAp0lORuEmPARkaDYVIU0zNV
ge85mByRXAT2Xdht/utwk8ugAP5Wtpg6lNIJi+yhteqkj3Xf+YSGFyqeTcWj22Yeysf64NXH7YQU
E7jht6+n8xbfIGCJbjyvJMBjrnnFlrev5kyEwFqF2pVTlCFtcGqzRvCYsHOukR7PjoBb0XYrQH6I
uC3qn6xt5CV+V6qnmySGH6gmyaa9+0DUqh8upesNtt4UI02TiqHeqfUzwZSO9zsfFLJdkqEqdSd1
qaApsOtOmSJNouIPURic/U1HRVv5ZNVIJYYzpXHbVOJRMaTFPuVtZMsXMJesETjzts/5rlm7MTN+
OXC3Q2Zz3jKviYo8TylkwtSstLo9ppzTgqaYkTgtJnGy6H2fWPeV2RO61lqCv3IK/PK2zLTRs3Wu
8pFMvu7NLsaExv5Bjx2mIQnIOXGRh2AST1pj2rLYD77DCBtWGECCLwkb6RcjfWEDyxwRHx473iu4
Rlh2EecE0EH5W7kIpoQNotjCYKehzxi13GFQNirrcCq9FTpeGEhmeOelGE1tmqfG7vRyGU4npoAj
Tixr1HW5O+RlsRZwV/mHj6KDs42qkliBWBDxmc4fMAGN8ptBHtIlaxzTznzPJHIsxdkC1q2qwhwU
TyqzDBFR19NKlyjmQdtdet2BbSEDsQI0MhCFdwGb3G16c208n2gRYpsU+hIio0BXlhT4/bnob3qS
YCqOQd5I2NpQELbx1Slrk12dKSb1z0rNs4kPqiIo8VglYbH3A8nEeoOfJnfqf9p961b6ocflcp8t
/Ow2+AoUS4kHWahvstdgHCzKks9nbPNBMwQ3wsVSad4t4NY4CWp8Qr3A8/AKoxBnsX160NSQrD4P
vf4Q3amj96daEdbL/N41592za6ui4RfveClfWATncttmlA1HnvzsFybr2AFnZYoPzKWGACjhWL4+
ZyNBNrbEOwQ01Kz1EGkzKusgOLkvtWzcqNu08/TqENGwmw7HYLQ9xEjVRvzkdSl5aBN6iKEoKy2A
3oyBSU2XYnAJHOinpDSHbIL/DvQSp5wvKVcK06Rvo9UTf6ialH0DhEZxCccI/JTv+MXJpLPv1DEb
Pr6DFEAN0L/cjNIcVDI/2+kTGIznTHgONJUWQAYAD6Z0DRPf0Q1a/PTFDxdHFhZrlLwTxY/cL5dW
yUpEKWGC/YFD9V3D4XDTX9YfTbJjIKQRaJ/8GROqrl+JwG76NX2oqCngcKa/Gogtk0UkeVc/gQw7
6R4zwVmgV5ay/7TUVDqzxGCZ9gZh5+KGMwcLXGc3SDKoABnXNvEbcW4RrVqUyMUJzwcbIJ+k12wO
I5hRRLR+jhX6oxgVmh24tgaoi485M1wTewbaumVQ+b14NJ+6E/d57l6akLB1Ov+wfx3CHXg5GaY/
clndG/UU7EraAyQCtcLUBz0r9QnqaYx1QC3kqvr4O1+Cdlps4KEXz3QX7m0GHhqgWTudjmdtZc6R
rXT9LVHW3U92rU1hNEnF5mlH2oVSZWPnB0uSKls19CwZMfasIQPOHD9GMhPqzItKPHrs8o3SNULE
h1zjdJ+m2518JKjCxE4QDp3l55Xtxwre0o7xG5C1kHZM6dKxr8IOjSWNaadm3jhxP+MQrwpwFizX
LkW27H5i7PZcpLIDhng3kIvnJVl137dgZ+LxMrO1J0A6YGtr/YQMBHOqJ0P79H9I6HTK4wRuMJSP
DQLTaJEh7mZfelg++fJGfsoobSMyecYfCCNvOpbyJe/e/O+buJfvpzLNcQTXLNWmdFG9mkqIOZ0R
yaz9VWapLbUHNmKBYmGEbXfta2lHjeSR1i3zWrsxMKflO1908MSc7JE7nJwfGj1WQ+mMm5wDIvpo
D69b8oe06txwijg2Au642hjTJUovtWR5MtQfzlOcWZOpdAwl/4levQagZE/YyA+bzRYDBpboqmw+
8U/o4D0tje7jD5PxAAkOaQSpQ17MnXOMAxP0IKDiU29asApvwVMEc/Iqf6xIOtkVybXGjkdUIeI2
o0NjQ4GfKIOK1aYgGrnt6/rVhPlfeSzbxqGiNDA5SxHdxwVgRFsSVuorPMxflPuZSe3XJBEKmMBq
i7bv+oicl0eHRk8sC92CF1Kf1lCAuNwg/U83G4y+sR1PHiL/7nilNEMly4ZYhbvIBLUevGb0hHjl
2LyAb+JHJGGC0BI1PsB2oYMhGh0Rph1xXdBLX4wo5CuZaLSHBI2cH0BYQvA50VYaUPIV73VerYU1
LYi3MCk+8Gui+tHpQUNZIcbhx/Vnn4ufSkfNnzGJhVJpliDo31u+FsqpXX1h3IcnGsxba0M4dSGh
MqOQGnU5lZhS0azglthlBO0flVGXaEkY1QuXUFMO9vbFh+raYP+4ujDjUbtU0+r6zrRT9j3L93ch
cr6AN2A9/NoaPl6UyWobLsiqnWy8NpIjNswKWjO0ShpZZOh+xDM4Btg5WwFsNz1m8vaYwlW9QB5x
Noesgq3p+eoAHHPtjqMBeHJe/VgaAhLoGYKC66FElG+erOKCCVg9wsfKVmhCUuAcOWHLqRHVriue
/8is3bFY4lgr05EHPgc+qrdulK/e6UFy/xq0Uv7gCT0dCatLl+AtDhYgLqexHyBfWI1CZjOChpp3
hPRX9f36M6KZqpwCse3cLFBFAzqqP/NN0oCVp36Lfjghhof9GCFn/OZJPiGU3pveIHJi8q12Jn0u
ocex1ijkpdKUl7RITdepnMyYWtHWyvs2apu7lBiqfJKWh5yZrxKKB/U8432hZsxhl/lRvJWeyHP4
nV0P/Hn6FLcT+TjJQTTSpFtXQrUcXHO7wS+NJ27P4Ps+M5BJG+hcEeRQ51tTf4xVRq8IR4JLcdsf
IwLu2GTabGyHpGqdOd+o6eYSKjE079zQkFaABg2K24Ba8nPoEjARRY0zWAxgHCnfXZWigtP4sIlV
JaxiJQdJSO01d1O/p644zMMnPfvWW3QOLysoNswJVZZxK40GHFnNuwC8hnxIWaJeCc93Ag3RDR/r
Oef7+WNOPMupNPyll9XB3emXKuM/theIct6VO7dejAArskAJck3u3V8ffSL0RmYIbw6/1G8ImB1p
kA7t0Zen2/jU8Z3SD7HtCHYj3bhcCm39pOjxXVIFfbnRJdmqppKum11tIPAXpdlNb5Fg/3bdSSX/
RIUhCnPKLbTio+2XiyJkedcRBQD2cvYHi9uQRqw59OqYZryndGiNqcnIorZEEuFNTEfIeKPwuNVx
Dq/9xAn4pUOAJBoh1NKXTZs2Rbyh9WdxJjxCSm4oMtCxEc0XoWSCumwnJ92t71oeUaTTLX0oSbcW
1lVjTK4i0k8w1sWUs+MgSnTzimwyt+whLLeGoqJFpsdg0bidz/nYvf5rInUU+1vuJd3ln1lhu7/4
B+bLHxEOKhV6Q/IZec2moO4E3ZMhYXd4ydYUqsTDHG8cc61KufldFH9gYyLwoTDN3JzhLWLqxZvR
rl8QsuKKz60kNXfmPaLQuyWZquJ/8rupT9PK2+Jh6t0R0JK5QcuG+9avuUskOmMKVSL2Pggt8TkC
bOLM1nN16jed4UzM3WVHK3mA4GaiHJWQc2jXylDH//PqXszX3eVz6FaugKJ7anH2C1GdbjSF335t
amn2XRZpPUNM2Z3Jt7L4dFxzp9r/6UqL4PPkrBJA/QU03DOObrvN7xG0C/jTzI/zGHx0ZKEnOpoW
lnH80S+btIhuyfCta3oG18YPaxAqltmRZw05bZVn0b/tGeefmqCa7sdwwWBtwlGuoShM1n21iZHa
y/JmTYZT++Z6CgHHL7oTu3I2tuj/2j7l79AWpyvLOFmCwGweDND5CivlM9bxl3aqSNfhz3lCF9dC
HA0DFNN2VWRx4IKqdivhfP1gBSnmkxbhn7ZK0PMIMh6DHW2Z+4d0VHIdCh0wfFaWxfFGaBpK6RHY
YK74rQxlz0ck7a59fEImCAuAXAxPQqaHWzU4jeGtVrx8/dAO4Y4MYInc0tT9AdTRxYUNJKaAgoEZ
nQm5Lllu15N7NWPGtzetFejmhcWyQ5TxWZ/LKn6sOGzOcD8pq0GjwUdirk+sJtr9Xlswhnhy0IOV
VxLVmsJPHcuaMS0CEfJ/65LvqVIFMNoq//rE4Z/sPD4YeGDZecNFOw7tLQwqEswFk7LobCbsaZFY
INu3lTazQASXYjd2vwWXw6QQHUKd9UcrSD0HtcnRqREwJQ9xUNOX9qCRKiMGsZfa+A7QdHzUY9xO
Wpn8HzRisTP5vq4ZAbkbyOb5mIzbB8IGR958wqygNLCOPohah2LF6GkejtYlejw0A1vC+0XNX02G
oLAVOHhHj/HAbfHpcK3mjDG6/EesXruSgWiRQP7KEljmOuV+BILIX7UOW1tY/G9yn0XsXb91UFAn
BQwxBNkOw/R2ZuSwzuyCCTnSiIFOZhPur1T4tUiwiH9SLwHHtIBd46GtLCXbEuhr2Kq5lxl5PFGS
HwX0QJDUfhBXRHCRVnxCUvV2IuRxLb9h1NPYqniDpRrAN2AKI1r8uvbUN9zVXdG7F4uPiwB1ZWYB
mIBpYpYaSYbFcjqB4ygWYQAb8wnKwhSutvgOI6wHBuHyTKzxxTtA11D5n+qEWljMgAQz9H1RoO/G
5RsiD0ByRl2SWhSgG3fVH68g8BDkqhjwAkKWJJToTzHXIV/PdNF9SJXTxSb0i1wYgV3V7oOlQzoG
LUBtugSKw9KkJb8fdMVo8Di74/ebN23qSfr/Fqf0virHPmKHf60jDbEwSP4JlN1DgOvJ/i6DW1tf
SsQPgU/Ivn4lNVP8d8JpkVugidIetdXgoSQv2BjP92oZ662t1ZJ7faT4FNT68S+QRyplMkK0VIgQ
lRfftew7iFRqQ4n/YFOjdHD+wQM7nMy2u/XoTEjMgATT1+vJMhTK0MvCy1oD3un+wsD5YaujMCgK
/WxSfcS2RE2pVpDEMoPYozXc/wb1coaKI4yq+ZMUHRO4tF+eH6Y54Nos9Ribi85R8bFMIBsgERj1
it9Sdj4pbBQ5ie5hxfCSBhv4ZIZhDMw3XO9ldukaKrsOPw+JoCT9VcyMq5yhy8l09hoBDoQyy040
2c+C2A0LCFQVAa3Pm5G8iK5vcYLZCh/REHGeOheMCr8hXpQBN4iWVtuiXKyiJ+9M8BHP50fYzqVr
9YLRr7rg0Ig8dkpl9lryD0vjdM/qsYF4cC3xgqB0/KPCAnlk16Hhe/ECqGfBBRsGvdi5/797N9Jl
o3nZYpOYApbOP0fz8RGIk/K63Dm4/f4qpbt5StLJ81QLANQgq1AIvUJosXsYR7T5mbBYompHozUu
SG+tlg4wAbtPH4jocbdg4FfUR9i8TTkWmEU8q/FkOc55mLx7/fahEKpYWEn7r2ragjjPlhjlbgWl
Y5mIF24PZCZ/Kb1EdlLhhzPsu6HYSa+AdADJNZCu4KOV31+FDbkCtLuvZVolg9Pvky7ythz4G9p1
VfuEuFu/coDLTWZp3WMPmvhyGXO+wwCSucfJixov3kutAsKdbRhFLLvg/vHt11O/Bky7OuRZJ5vr
If3ifq4d6QcT7+j1ayWIpsVxbbm7sgNqga2VzBq5GOFGS5NjpQkTrfp548oOcVApxWg6YJmECas3
hERqDpEv8bhEUmxWAzUD5lMeMFtq3r7qTixxDdYs2nMeviWahsjFV42qZty4+KmzOpDsEGjtmX2R
QYjQujeylDMFzkSuRkKcqvvZ5YLguNb2/rHf6EhOujFLASCrLiVqprjJjr9RT7MeLL/aBal8Zd5h
DaFut4hS+ToLC3LHoK+JuqZUhTNPQauC9WIEe5qV6+aCm+rPUt3EirCcg0aDadBrEsz2dIQXCw77
oCwJtBAC7LW1t4H2YAe99rpnAAy+yr0FqjJe2rEtJK5ZGYYdUYlLPUcVvwoS90JLyAigFghWG0+u
QSj2mWWnXGHfFYz+WNosiSn9vqWrJqXN8UiEdoSiy/JMnjY7E/LbT7XRsTbKtjpKk+xx1kFKYjop
+pCDOzbboYCdRtjNRcGCVTAYpYautaN0gN5A9KBfcTCiKX1lpgAd22aFqEjgYSDNI8EBvXp/GhSi
Lakt895IZKSWP3kEgdmh/ruFEmN834e5bjSUBM6A4bMAaQG23tc6KUKXy7Kw+YFlOplaMoi9Yn5Z
MuvzZn6DIR229u3PVT2CGLtK3pr4QXunk0AsdcKd8DvQgM/tgG6DC+LLRyAFnZ8FfF98xFF3T/we
gIWS4MluJpKnFW59Q4i0XzIUe0he9cZRmzmM2+s5cZs/m/sqFJxd5YJgKHxAJt56ADOWVwd0qlCK
dxnyRqNaypJMmHweAQi5bSUK3H2r9mfOeEX6VC7j1Z0Iiatp1T5RK28KJHZ/uBLwnx5DVnOVqQ6S
82ilN4X1wKFK2G1F23+fIP5JfV5mWWPm+q5iSEoePxqpR9xbT1JueHWio4i23QaMxXb2K4eTRSki
EvSDN2qUnw2+kikfmSg+Pg9KCdcJByN/Z0ykhNQhrz28g3Ye55Wfur58HwDKuhxK3CUCSJqoyiuU
ElmCZhZUuvqCMD3imq4OjHCv6mrHp0WNtCZSCfhpZWHZk4S8tEROlATy4P+DXpKWacGwONymmvNz
G7gGMxOUGoeV8CbRkuI8iBC7wtQkr0XhLdeinhsy9OZaO/ZB8wGmKepTykidESOauIEwX057i/69
rhdHFrCGaTTs4Tn6uF/iu0SX3Hs/YWBDKik5IgvyA2KdklLTuAF3GheRCWHPSnX2rQf/VDKHwifq
fBFNit65D80Rfwn/ReqA7NnkxNgboRjYKBr8ApfjzJvWIt+A4bVz+fynbl9dtYW313e7ZDzr82vC
nPP4x9wpiOIP0y9/x0Y5adwMcvbg3sam0qZDcDYxXg5+g1p6TF+l82oOWth9ygCoq1StTbb1mVDt
+ee10xH0qLjvGrV8drjk+UT//J/jZ+q1k+JoMYfARnpSbz4jWSrBPmNmPtYL836hf1Dgsr6JJC2X
xV+jV3mYfyzc8ItywlysJGHma7/6JVwf4i9yjhljYSBOf3Q57vgsmOE3H88Ywt0JnEn/NKOyuGE8
vovEmhP2b46BLGqTeYYuT8oQk8c2LMzv3gbwO7p1dQj8xzPG9WQeYOLh18QlnhTMJXQMAA/6PXqK
cyIiO9T+wCbGkSFcNByQaCSN1hAVP504PkxiI+m6WGdEr0ST9W9Soqrt9cHY1HnJPUkDVLkSiHrW
vjWUJD69kcrirlIxG/2ZjrGO9OV/LiLd5g/pGcExc0oAGMFOO8C+LSatQ9y4VHzySIskIGgFwiZm
mH7mQSsEuM9omOEAzmfLLU4LYl1B1m0Ow8bbS20KHu1XxXvjpSl71dKpZ0VO2dbO4un4LzA2Gwsh
FTyO3jITYbjaqXl0GexrYgbv/QcEAcfHwX72dnWq5blUgpCr0iQhheNzCn5X+s8WWJVj7QtICldt
+SAP4W5SGDL7tFFGosOatmDMN6I3laIkxSZJknTNGXJ3EEAZdDu/7IwnoBltT5ThKVYAhFdfA1va
FDod0ShaaOlqYSahbaYxdA05H+RAKdtnSyoYX7bu/NB6L1NxEh4HK+64FvuMzNYsO8oVr/VWb51l
0kFgPepGEqtyeedv+is0VaJl/D4ARViXspV2M6XQhz/bgl8rPcyQSFvJC3fAfbT4Aeduv7enoghj
6Mlf8c9L8itdTd+wd/J1QQf/Du1MpEh69SSB8Kum58diOjtywaSaFi6BDeaJFhhjGxkft8zsV6Pj
A/nDBH2VVtMtn30nRWZ1gBEkSz0HSU+Xw7WNeF9xJIPkFK1cj94YeT+rMdqDxwBiOOFRK17NyEDc
fWx7Tc75jWaV9VLqo7ObUQB9vtcn7oH8aSsyn2ZUGrWSszbGMQrBYnAbdDEDsV0gIAPx+dytT81O
xXIaf9WaYAoHnJUAOAywdi4CbO8tIPaeldvoqZpU+TiSPL5NXxuC0uvQSlAfoAl65VKNg8pq8geW
xUGHbPgQ6VwAJviXW6qyERv4XfCBLrUoSuk96fys5Fj24cnYWh+VoifaGGWlacqlVFQ70GEhJ+Nu
xCPQA60CNPaYpCp1U8d1J2RH20ro6ho6xCwc7LtUEzNFyoPzqXiaJszbnyR4cRzQUekG2jh6x+ai
SMbA4NeFBvjnOiCp8ZyyX7SGDh7O6cCNeCqY59zZ8cn4AqS9JTH/SLE1xtAQ4+LiQ4Pd2t/Xr/0X
11p+uLGAkouHltbiyxU4eKwq9CTj6jJ/vzNG+sGt0Q3WgUNe3UKMqqcu7swhCqBY7eXDGKqNlsyf
aV688LwHbCGkANnNwiN7VDmqGh8yNgtIOLxA1k1IPj3X/djfDqBzHabX/yjU4COAt3KWMqnc3fr4
ksPd6gsfdxSjM6m21IHHi/0LYVutdRyX9dUtiMTAmovb+OiRePb69kl15JlApfuiq9FzoM/Sx0ax
iVTz0aVXYRe2G8RlJYrBm/hMndf3DPQQzbfulkhKhHpzNE7NmEs9qu5+8LMp4Dm3qATHxp2+cUAN
yrGZ3UxNQ9MTrcLoRHHacbje89qIg40f+b5l8AlCQmqxW21l8PRAVLjkJvhToodMBX24nGt2StJS
4FH9a5ctLwaXwtfATvpem+m6tKRe7ICFz0xvEWav/QWHh2RDw4geqxku+iTKeBCFvpL7wuT0f0Aq
R1swjtSSDAieS49M6LPtHADK/pzLJIENp0pAHBXPV8YKYLM2l1jfHPP3EXiR3HiRlz83yfpGlOTa
ETsj3teqh2dBFtt5Q2D7lTGepTUfP1ZPX6lH16lmb3+8L86xOrLknUBzz8XoM3eDlXM2YVhmygXI
Csyr9v9mavRokMwzXw5NqHeSAG3iqXMN8ts5ZyvWZ0s2Ws8pbiZFy1rp4Hr3iPAznypdRw9KDgRg
5c28CigsQYF3c62dOcIV590c4ql2etxe/rd0xf8n03wwc8+bWT0d9/RyrJBDfIi6d+lt5JwezO49
upkCSkYWHqFSLM9PdzDzPIUgbjYqfXtdh8G1UfJfgSrVdxvSquY+Z9231+uRScJnw5wADBtApybt
aZawfv6N2r1AI4w2TpU9fn50nBLHndiQtHB54R2AKMg1KxPmgmX5xfUyatlHgvk1k9D+jubuo4xb
crKJIGJ3pxPz+n2JmrGymUPIwsuk1Wa6V+FJ2Z4iGGcCa2z3b4tSR1tRx61OvDuKjDRWI1PB06qd
WV2oLnBUS+JUPchhUZRyOQ97cSbnRtb00Pk/1suOLW+H91vrW/4JkdDCHX5kWZW3DgBHQ6hYpySn
lSkwsimAtxOGa+iZx7PdNQYB+RQ7SfRE2XJuMPM1EpOMSah+FVKmQw1U8Q7K81t9kRXklr+G1koJ
Hg9WnOemjXsZ9k/Q/S72kDCHbzqtJmKDE7isSizsITP5Vr1hDvRyVrbNjWLrFs3upGxoscg+iZkF
KlqLOgsirbENfUCUrejTF60YwEt3a0Yf+GpOhi/SaMBCysrDK0jBn4BSe9k9cDfVtjWRFl0VzStn
RmGY0Tj9dxJmxiPer0e5omZxc0e/1l4GAKFFSQqmlonEp0jMAyv7P7vIrSXBxCKgwgXvaLjUhQwT
aTI1L5FhcnlftiihWVe5L0jOPDCQJd439z+XZL/FKH623I0/ELJbiFmEScdlSXk5cvGkz7bz/eMe
Qj8tLhTQZksORKYiiajPunuBYxwO+koRXgOWXDfUrs2M4X7i2JVx1l3IowlnWp1mKis0TkpE9vh0
7nUigdb8SXzsWltviv3NXT+bgxIsy2B1wTPs+ZL8FBYqBcDplKucg6kPSQmtJLE4hlk2kB6rckdZ
4yp1Iv+uJslL4tuDeZpuqZQfnxR+6AcpS/hX3uePUz3oI6h0lM2w8ndm66vHenC4aPJuEE6Al4ij
LeqE8agxFueUv1BEzqmgelFetAwcPwwLGAHMuZEi/K/TTM2nCpzLX/ulw7JzVWpcitgXh3Czf3ec
ioM94tZ8K6VRJC4ntfOtkOL6DAlicDWiA/5eeE2qwiwfF+tL4xC15hfKDYouJcpUAtKXDRPUmuxy
b1En13svYkN1/cQeF2S1E5ixXZgSl0iSDcQVOMQgkJe/SJZyZazeAD3PKXeaI+Zs/icG9zmkoaIc
uZZ/E8xwrpG7bkBFdopL8vhds4Le4odjl8sR0lXFlEC/TJthsPtPq4ha6P8MrSbnE+Y30KRjMju1
zabC85NjXBkackHXtdRDjNdyebFVPKxAgmz8Mfh9HzYFHhv8CS6A1jhy2wp2zE7MiIdeG+p9iXWt
HjvrEY6ncD+lZ30CZGslSjEqS3CtpN1oPxap48Wpic2MfY5PSCozq8084mt9aFdEasg34rQ1yyU/
E7wu4ajTH7/MeJJ55pLOGe5SHIi75JoIzF/w0q6RaGEAnKmIUnYZr4NLzPnfUeZuSsTmOKbRT9Rk
05NOdYRUIZXqRzp5/gRbnYLf8gLjcyRm838MC28kook5cSvdouqAHKIKVM1E1K2ZsCdZugLkVWVQ
rYXn+NHDzQbhvIX2GvW3LG5fJS9zZ83Be4PbcbHKceTjrnlKMh/r6MOrJ7mLkEsKd2kvQbts6Zi6
uqIjMcT3k0f6Oi7FhnZG0qpCjNF0CFqdJT+FdLkxBao9SF2RCpqaxOPhklYh6W/pZx+W/IXg8jNE
6QvmygkRBfZ3mZMsKpnuZb2iNR+YnZgCkiXcbGXRirseHwU9AoApjp5/HS1fdlssOL1wGnJ7JovO
StS6axva0TNF8Kz1xQ4YESdtqUNqxqAT6Zci+Kt5JKWriypCYW15ZcEdsdVmQXNR4daDZMdFSSC8
2VNBcZxAhC+mVcb0wmtWWnOPuq8E8Y84pT7wLcHLyqEX5BSXThvoVmd2TSfKbvgydJ05QDc1PoVX
sCdzvI0FITDox+MY1Mmm5DHuHQPMPJKe8YgEix9NQktIEEl2Ds9OyykzAiBAzT5QN1007r56Gwrm
WIfDFOtrXcbalL/24MH862yB8pxhg7lf5T03OPjrumjO6b8iFisLNu3WZ5DN82NRYPbbOUP3jMan
9pzYfRKDcLi5fKy2Xqv61Kw1a3LnIoHYZdhDBpNfVCnp8hu10Kjmyifx7xVaE2CAk4auB/U+0VOw
P3sLFKQD7izOJTQX2RCgZBY/e6Lh+pGO0xA+d7rBLVu247LGk2eC80BjNRphWvwOnf+nyv08agxO
Eew1ayE5DgcTe+lcFioH8HitDEhCCd9sh5BNGRR/iM+oGY/AggxkO6+faIlGUeIq32V5PX3SGbc0
+hRAgGZHk1RGFE/WONzQDn8CqSeI2GfK4Rnq8rUqDwESSNsGvYo6qktY6xzzTQuKZh5bUO/svB4c
3hLBlYOp80Y7dMo5O3QUvkbAPwDGUe3LglfgG2/ZB3TeZrfxxbFHrGJTRIMJGv/1TRP5QVSGt+RK
88mCuG/UGdmkWigdEZnAj9AOLJ5i6z54lK0v1v3KAsoE+M7WU5YaJot0Hf/nb15fETx8gYiO0ToW
ghvOZv+xsE5OJ9o7L6dynv/7szSSgyMtrO7nGGQrse2QTjfXCq6zQNCd4RQiO/nCeieFcI9BuoB8
/QYi1xSMR42NMTwnqWOYpUDoxmxfEav51jKDbDPQ4rrAQqaYvOBrfOrpzZhGyZp7Wvf7EjzkNgbE
nzg5hGaQLwSE0k3l17EoaaVkd1AQpDp3R8SfVU9/V0TG057cogN6n038L2I9xuieJTV1T368Qc6B
4L16PrsBOzZYwVT/fv9iOf010retDGrSqEYpwIMAHvXVJICLd8qUE0rW3l51aadgWlGJyc0nxh3+
402cH21mKK/JSg5pvPDKkxbyvIMZg3KdZX0rNLYXHctc2669pXI2MV/ynZrJXL4q//JO3VxGmm6L
NmfIbxCLLz4HSaZ9bY1UDvlXYRC59IN3rmiPx+L9to3aVEMMr5xclgXrivPoWLHMhhpYNotxL2gg
REzwsUMsgOkU390vMpZtAQCcsgoYfAPLJlK0rUreUD0fR81Ib2RwmNCic3nBj1IUef9U/OFcJ0fn
QyTKmtm3GvES60wST3M9IHHGjUgU3b/LPkNEETW/8RzYB27JnOwAgiVhjsFt6CHkTmzYc+Wmnt/h
/WC7IyLw/yBjb49Rbyu0jHui5rPjZfw6eImAyKuYEttgzB++FnuUClAeHrYCn/lbQhQu5iqRyv/g
ev1304Ie1EslD8o0FQBKjuNpLutRR3GtUhg9mnPpDTGO+8UXk4gkkezMJ+jeBsLBwYOO2U1+BV42
tBcIdL6Fw54xPE201Tmtf2aBx8EWYhDBc4TGe8SslqfPiGTXeqXWefKif3F2FsdnmAAYgmJsFFFB
ottxpCRnh1QJTscoYu4/mwcV5Ji4vL2p+0yGnyDKcNwjGO624UJ9+BQ6l+uasav6RQW6l5rL4ZUZ
wZZX1NWJADDr8hlZ8IqG7IVFClYKMZWpUPEXKdBUVY5Z0DTtJj89xg5GyPCs6B49c6iav7O1WQLD
py5xFfXAi3qbvqAixd3w2LPhxiHffYN7/+snJV8Z0fhNIBEdTC3BUiEPFMwnhOmcin0CpWOR7HO5
8cpwxhjbwoU/52K6K3rSMZRhUFpoF5HVeHq8TNHieuOKM03LDq7UliTYP4OBrzwa0lceC0SboZMj
i7E2uJ4aV4MyNp9rRINiKsS0ETWfnLwGSrV/o201Ru6oWNr7psTX7T0BtxKLsil7U5NNFgsympMt
WgmVjtYmIW5FgZJa6wizF/cdL/QPur57o5O+BWiN9UWbuh0y7gliQCk82BmvBD3saHiTLV0xYGYC
zK/PV2ce1Ob49/DRtxjV7tEsx8RwQc/hpMnT7YmBBB9BKNBGDuuCE42zsQekemEhqmnVA/zp3hH6
MJoqUwwafzBn1UafB/uDNON364dBoi4/H8I2c48Im71da7bopHujCB5rPROCdXUguEq7F5vXSu87
ddORtj4hRIfcCS/CGXBt93bH01pjji+PkDxOiuF4mmeR2eBFt4fXa7z50VhWz9Jqez/LROYNROSF
9ndXRK/Vv0qPXgc9KCIObJbWMcwh0TzM4mDJxWoyLR1zHhKaA7HiAecFH3xe6I/osX8AE8DkSu96
cnfeYF84Nao7nT4ugiUAjKxPPiH30XY/xwTjQZQjV+YdM/6ejaFGX33QX6I85bbjsc2xNyH16P8a
X7lluimqaMuird392FqP9HNR+4VqeCgNGld4xV3+/2DggbLHO+RZj6qLoZAgeNvPWBUMR2wz9094
44E19eBA8GGC592QTgWea+BZiMGe809AhyzBwdRrE0h9J6oDCYR+uQX7gR3jlojh44lE5O59efuF
oRvMw0XukVl1Q96qJoWwReAUDPkhbzTJ95goJTx1TLwl80srMEy2Ayzx2PWbo2klZB6j+D1DFKFZ
TUDRACA7xRiIE3r8lwD5B8DZ5RKpK+x2cOyusCfimnntBAQxx1Xzhh1KbF1CInCMRHdMbCc7kWiM
10yLb+mS8mghbgF34rI5zeGVtMoPtUmkfJSyOXRgByNUpmlE5xDgY+arpiIHFdJCH2lEyYlg4I0y
IjC9j3o90FO1xS5vwUmul9vnd38UPp0Jyl/F9yGuGS7IHdqJvXSJizEVGebl1aYNGEYjnE+B9m2v
qGmftVq9OCSw16sw3nfmvlG7Oobm1vhtHZkPNiqkHIrMqhYVXCvQDfEc7naIkQk/cL5kKXRfANnR
1kLmGquBSX20ozFe0gvHUagk7eI0ww81IHzpW0okAGWMy18kDwq9khVfyRDr2ICB+pUmYBVZ09cv
SRrre/zr69ps+MeMITpjN5juT99q/LeWRXlPsp7C5vmtXbSDskOlKB8jfBLl1gUF1UGaAk2l5yXl
zHvvQd7pKL+tQ0JdUwXhvkCV+XAhnSf6dhsCTxGVxqRwVY2VIGjbo94p/S5YvrEK7dbZ6IH+EQGl
pbQAT8v1oohnnmpd+sPeXM34GyseuM50qDfZQ4j6aBWhkCbY5SHKUSphxV9nJzrcddZhD2YrDu6f
LB9fnxUAs9zm9DRRf6UP0uSL7GqJhn2REvrhD49sR/vsnsmfj7alEADEWSdapSwNkp5xKxRFK8wd
38rvE5MS33Kf6VHq2f5txFiNMTTSINT1x8NTslcgeNnVjcvJto17m9Xfiu5inq/22oYY0gDZnMuN
Oy4ol2HxFWpfFavs8SH/i7GRo8BQQS8l6BAZlkIPVDGQwIGG1VshqBdm1kDb39izTKEbVRyY0WST
QF/LwMPUDOcHL5Rzq/obkLrPiFCi2IEonww+ivMtVaLBQInvFo/2K4r32KSvlBwdaOMx8835kosa
o4eQj4DWKIoFDJHqOpymwtd8NdGOIUL5e8VtsFx99KiLa9uqi2PUlfQLel020ljHerVBanJ+1lXf
TH4jcBMlhYuHo88pnAN1NzCH8N/hzxAZttO5vdkT2U7f6Fan5stUamb/o26paGOBNdJr2egkieoa
xv5rWhjl/aP+CWbCOE6e3hoOwnO7tImk+RBZXAUGhz4pMOYO7YPGufYO2jm8ICZTSGs62Ki5Kcn2
7omLn1YTo3Mj0nKE/VdVLzTcYOLNurOhpN7znszbG2zyI8G9vFAD+/99CKToea2NMR7gBZpaRj8k
ovf30LZNUHHQzlLmM9AAtMBQK/GVe0Ts5/AnDPi8Sjfc6U+goKbLjQkgvaqs867IpOykhV5kGyik
NfKQoFUk/86irHwV7SQ7N2hBi30ioHmH+Ew8O/3o2ih4CnsShygm+tsVBo1H8kGsqmQmN2YwJrnm
S5kJ95rN4LwNTnxryAAwvOlt1TvjFFZxeCwbJa+nDdO/gdoPv1QCm0nlYth05PY83RWV3qVbjO/u
LldKijRwRMaYOVX35BA65xBOkVInJnd3YBOwF2juoFSpwduATRI2F7UITrlDFBD3rZjBJpDoxC1H
OGlE8uMQ+zTErp4/9ySelWObP/PrlhREn8Z/DhLsa0fhvGGfYi8eQueYxa+mTrkaA0OsMbApeGdf
tErDYekT+OFg3IArmKFXvje5GUZZqEc75RWHxMNtFUBiTOUikQ8W1OQOv3SlpCfdJ8prvSJotL+C
kap/Tuf3BH6IbdlYw1AdOJTPgmAWRTS1BTfxp+g41Czbm6AOmBnK8BKlftnPpmasHnJb4ylpZrGK
vm9mEzAmIvJeSkyH7F3aEajSvAxFEtcnyQ6E9oADteHG9iRKcolkOAPTxHuh1Xh+jD5pSDBXOwLi
KdIP5ItGAURdcACSsQenMQowjmj0Oz3yAIQaAmcWjmHkl6kvw0kunROuy1ibvkFv7sOQpRbB17sH
ZxKPgikc8TNEg8YDHZJ/+XkXbj9TcsnD5zJlwn4YuWckcqwqr+ZUMucBtK4lNFphpMmcfRAkLjOZ
Xsq8EXXN3ZpwFlLW//epSnU+aaSyoe6xUUm1zVm9pZeyrLvcn9UCrLFCVJiO1CGptEj4e50daonp
BuNTSuNP7LCBY7q40weKwjuD4eqo8h5S/B2qoHICeZIwS/+XfGuIpnZ1/Z/CGglWZ+mVVBTrIo92
0fCBBgmIwEfhybM1Uty9jb/SHUD8cCTktHlzfKaiF1DqWfnYPANq775aXOFZtjGjd8maNPF1yOZF
n/+a9Y5o36HsIrEeB2WY+gQa/xh8o6QyIRU51PCsaWCNGSSyXrNwRxJFsMhNoO/SRTxcZwu1ZFXQ
uTneAxUEtnjShQKuHD7kk86lSzwsIfuf4GTjcT1b5XR2x1d4b5O8aq0bfrGyTKPmWz4LvWLQ8weZ
RrE1f/3JiR874kxGuxhB+fXYWWkNgSB+5R02vTRZXq8jG6Mnumy+C0EFLW6LZO1WeD+Fiz+qv866
YnaMljakeZki4ss5k61j7E8pGlkSdNYY3oYss9db4+gb+EIX9mI2Poxvuw6Bm3vBf+eZZOJLI2FI
XCMt8Ui94sgq65oVRX40/wWMrXRmHzE300/vYyAgAoD+MoIbfguBpxZg1f4l1nihZhY0VKKG/g7e
AmXiBHHLYSvWJ+691mPWwXNH2VXdfwAFvBymVhGH79xH3d1KYcUHyIZSdichb1C26g3u5+a+758v
hGleEo92nvaXV2jtaL+AI99ejwIZtb249peVRUdh1jQptKMmOtBKtDezs1aJ5ubXJJH5avfx7mLT
akRGi4uBz4Rl2EgH0l3TLkfmXYq0RjivgiVZRveDd8o4NvZQ3aGlVqv57e9CuWsn2ImbINQ6Bwl8
EXAy548qDyFj0hbSMCUnmgenUzFyaOdp/F3785NM1id7xpEi3HYuaGlo2RclGXCq+4/V0+y2cD1O
3zCFVixNUjWya+kkSqGBD/nKU6oy+fDW6azn4mfKv28IsksbEKtwHwnTi2YQK5DET4mMBEiIV0xM
S5TIf0YLhumBZ5lx1Vdb1JjA4vD0Q20fpLeWiWWNcpXLF9sigPDQHwnUcelkzw+t+RgPfhRGiA4s
ET+B3uSimZ85x0sJcuwARGqlG8Jf2O0Sd5cY/k+0WN+m5ReZTGN/SQPj4fGLpV8fF0T14vy+Eod6
IWW3eWZGL0srOPuhAJdusUg91gUS5Ih4MLswuVnc9gtd2T+j4+umsD7yQn/RB8nhBHPB0GJxGs6e
7Ylcjany3SIM57kvWCdiogQolyG+tYAworzVGZ+V3Y6fLNKM5MNQ+awwfF/i2QdS2PGE0JIHZUF8
5MM8a9ZKhBOqKLNOWZMG66rq9iNCivFEeNNmlCWO0zzcWdMJnF+vWy9AeYTMWVZjYQ3l3ZjsdnPW
QYar1S0Uh8xXWsqjmYuY5FqqdKUMr0xRfmQBlHcxO0Rl9sDDLu52UX5cw1s52RVPkSqdzt+x0MBL
35qg83rEJfhvIA2kZd1+KZQ4B8cmtHgiXHKjuQZI4BvBm4YRVTOFCjIIL3gVuGnXxhxOIBoLU9vV
Fc2XsV7Wxdlw94XRHB2v5orvmwOMUe8f5e26bECNAzb7Y2cwSfxsvT1eEXueK6FKzAKMqVBg0rCg
8m9jp4vhlJuF19hJBJ0/eyvFomrM6zN2oWL77ov+cRM2VvCikThs4oiFrix/tjuXbdTMDRfV/Ir7
o0qInJVnKiUJZyqpiUH+XKdSJWrubTNYKOXb+n/+oUQL3VrKutYrxw2EHevFQMVqwgflgUHNa8z0
hfRIP17RPdsepHh5sJf1Auam0oJVTSZrgHY3arGk240gW1dbvQlRMLDAOR7U/Q0BUWpVT1+j7c4e
0Phm+H+V/8olcRKcdyrNA/499kiRgzHJljacpa4+cfp3plEWWgbO7pSfyvlYS+Ng/F9HsV1VoWLm
1wggx6CSI36bsSspBYEAn5sYD3KyLnXUrS6E4tNeLjIZVueR5LD+uAM2j4jdd7Ni+ypoQSoFu0fm
pwf4wQMqFKauKZd6hdMnXsY5vYDjXgG2Og9yenOh61DGFuhK382C5a+6j97MTo2mLtVym4mY15RU
r78eUEkODS8OlZgaJOysfQMzMqm1BFI/1RSx2Zw+HvMSuvgIQRGPFsFF+B2+VfuCDtgDKxmZyunY
ihwbnXsS88jxwPZP7qTuqWSvhrueilIb6veloYBulnQ9gI9oaRn/iigil5cUJhOQRyDeL3yQDdhG
dL67HKuc3h9raXwTwbNOs7j/ZiCpTRY8hhZTtZa8JNQbmekoIqVA95xVJnWeGDwKtK3B9qgLBQOP
JPoRVo/HNFNdPX47ZY3x+ntUSM1ejEcuTMKSvbNKQ1qEbLFnAdEuY6vLes7pD+Ouf2GYuyh/YEPh
ou0f9V8P0ZZaFRv1b6DOWaGLEiUyfJIzA22HtStr0YtgiNIeQiDZq8ddGTQtMXyxhnv5MmyXc21v
KWBGcfSzTf3IwXr4GFbXlhbaMzl9yIqYxyWjplZjMNv9wP8s5UPEaqeo2DCbYizMgHyOS0sPnV6b
MQQcnmNc+hatF5yV5nAXwhhqSeSeLD3EoePCD9Ngo00YnQZBhfQ9+HUnRzbcX7r0sZEsGmWzoU/9
HvqnImBc/6qEVnH2aZJgDpFWbwvwigMpm1ej/M5Kcf+6Epi2g/QoauevnHuq4Dyc0Wj+YCxEI1Rs
a7vLzLrWwdkFqpyII1YZec99GJnzVMvvjnJvIkUbLrdrniD2lIBV1wqhwC6JBe+EVCSkEajSpV3S
Rlm1L5EDT4p/8OWq5mwfuLXNtuyL7QocBzC34mGaHwtfM79lIpizYcHSEEEKpXOVAo7vNtbPt+aX
pVgqJRZdxcf098Qi31hOUNGPLJlBJvRANXBMB/v4ic8i/XQ3704rr+59gTFWTXlhIsGgGMJbUKcN
yMjz9xqiCR8rUX0orf0hamDIaWEtm4hQKlkUVJuS6mypsDCuqiH3XXTmFeJwMfejOdkUc6JzeQmY
t+oD2VpArUhOvE6PFn1AuXjbG1zZPS4jOY5TgoPm12lqK9y5SOADshPAFDPk3mLvpFjQcec0Jwgp
mo5GyMawa8drJ4LkF5g4+9L3p/iDjbczP9XE9kb0rEHFACQSyfMrCtw4QI54aS3paW5wXWeHhdi9
VubIOitHRYsfDzR4zT+m80za6SFn5Qe3aSAlR5G27yPJYrtYz5NpDVamCd8vwbYWEI0kaRJeeFJM
3sUBfZCcD9l8K2JCQdFsXbhZZzwbypKYKjSV31QxrHV67AwaV91UPr+HsFFL7+Iiqc8zWMoIxGTM
6xS4h2NqN9c1eiknrccM0TLXNUqZuAfPqU6dgLNZq5NkJHh7m0VHT90K5j+HaqF+/sYarBFAZNCD
cjkBP/SL4xTMgVa1NCCD47ZjWfSZsBIQbEhkZ8zUfcXabSF2DpDWcMQ8bZAXhRNGMAo/h7PGZ2qD
q5n6BKJZMWxxyzZcyg/b4yAvWvNfqEp+b561tWcRJd0LOfbBYzcyzIt3jvVlIGAKZoPg8892hU0M
rTuWY4V+vgYNy+/qHYPuovUJJmV0Q8Ic3AJTkIMZLeZVvtW2vGvUm3pjzcHVSu7PBYkvUDCRItAQ
8+TQm1PYkwy7SBksaZfGo99XdFWLGfDvpNbULUH7zZrzEGEkvfQzvlGfJLDp0LXhOzv4ySY3ss+q
kNrblblCXR3BCUk/5v2gSXp3xsj9dA//PyGQWiZcwyOP8lxesIR5hKOVkQ9h7Y+9I5xpXyX0t5gs
gTO82WvF1+z28OPorYGuMA7DbbcVj/a0ehImEyS9xzpy5wMZzoVrrsWJipTcjwN0wM21U9g3AvIm
6nmoGpQBxyWcrzehyqL0jhopcdNQGOSexRxTa0GTBgATOvvwWlEv4PXXZBMpj5beovugcnqxclFV
aKi/aXLQL9L+J716MIlCsAoQk6A8E29RSS0ylQAAMMmzVP8PBZJRpZ5uIq78DKP5PCRiH3m0Sze8
ajfUYdrIrDpaxb2uI4SSGT0gkhQYjO/ZMYuPWoH9FPzY+HkO6PMOrNyIFr2+c0rnGbxkn1LluZSm
maPVuHEj0wwUTBZlalORqd+8qsAXNiXZ9fmocJ9WwUXXwTOw/jAQfun64dAA1Co5yk3ziUDU3XTq
y8OXDhcxLOPxfpD9rWmpP+sRTJoM2xslFD021egjpseT8oLmNWyxJPiiVeFScWgcnZlBx4D5xBeV
P3wJWSzJ7L8joSglrGsGU6a8Y1lnB5HJRkJ74eLallY8gjMNFDLAFqgNE5fc87QNC9XxvPR7a2k7
nzgpSmCHOy6iMWy0vmyh16zw8NqY5LutPpcST1DDXSB97Ca020JvZNoSG5fEU0kMByP1vZ/foYwI
rhqhw0EwQRcavLzSDJW0d8/dxE0sbYkMoqX5fSDg11AzKBA6VFnKhx0WmsgdqRoI+4LsAc4KTnRC
eW+EpZ47sgD5XjZp3CSh8a2qcs6PorMkvw+RJ8bk4uXbrGz06gHHpIEQZVcufjt7M9J6KWMmd6WM
8JQ5WDbdFvkJL8kyxrE40Wv33cqnRidpDCWhOzWkA+nuNCH5a0Je6lL0d0MOrPf6RIry4ZKfpQ0C
xDMdQTNuE45ZsB2nGECieKdH0cb1KYtByUmiGByn6trhAmJ/OC5YdLnqc+9M8VF6wppyZiGUoXGl
va45zvlS/mg5C3E2LqYb31Wn1wFEUGMacOrtNwa2IBUKoZKbJL6kq30+nQeR65YqAC+J7kMG4Odw
rOXwk0DO4IncUe5If1C1ZSY0c7RN9Nyjfd78T2UF+9gVcwYRmQUTGwrzqJhzlgxo9UwCSV7MaF97
9icU3JfrOLNJaLIsQHBsVrbXUHM40XBk6cMGDQ7wAUHosG7Di98QEkNIkyDay8J2vShO9GoNewY5
if6vYkJNJJ9N2BIgzfooSVKP7qhRi0GnFQk7V+AtomV8GIw9+EvseXsjzXoOhuvCv+Gzu4xqjjsu
t0W08ZP1o1IYRNnOJr5qveKqPxxmpppDdY3vC1B+nvucpAJNMMLRwzXqAfn2aDy0dRKkZrqD/hcS
nwF7/SP0L73NqYdLzlc+u2u0VSv0cWTFf0PlxC/89A05ThwS0yA50tnBiCNL5flvx1xNJzYQ5DLt
AqFGdde9IqdS42G26Z0azWukcIgEmg1f/BhiKF7db04Bz28zL4lKeXZbmT3wOtTui94GZok0oKzT
eFFhFOYNE4JWtQpfZQxWXhQOCXL+02Ml2riR5I5mzIy5PsGruwlLMz94ppX81Z/rUmc8KHa34Lkb
2AQia2SQszyr+HSLab5WHHY5FgiY+81DbUvC6v8A/A/+N2xaG5WqsnJQbwjZYvz9hg67Z4sNppRt
dYDF6dIsPdKMDDMBhz3ve28adFxua5mTxqk261t9NPeKQKoZnIeIAnCWnx3qtjbwmTGErRLqn2Xf
nIbwzuO2A7+eTHDSQOsZ4p0nPcaXY21f65keo4S9gH++2YFbi59o2wgkPUC/flrlW30oKuUSoRJf
Qka/AQO9oGqGmI7uGWOIV2CvUXTTneeD+KLb7ln+COYenAbU4fITDWVBNDUUakR/wraQi6WNZFj6
ZUiPCaU4Rhgd+6SqRGSH7AhIIkrwJEi4mLVeoxV3KEFTVX2ckOablskIH7mnDbW0gv6wbavl1kPj
Kw0/jH9QjYNpNX8/b/tpsO31xg8AUdJW0osJ/Cmdk6/RNXX0p3RfnVteqkrXzeoed9FbWpRwaDWS
NL7XRaOSKYz0YQ0sIZdxTrf/gBp9y6UmXL5mAhapPlsnQ4CjdqyOXOiUS6D5X1pGR/ggUf7FcJ7p
itDZQ8/+88R6qmY1lvSiz9Eg0lqNu2hYKkbmIb0HifUnThtgHAizHBpw/pez2SrBU8Yorh/h1z/d
1Ic7Cj6sMuYZ5XbpghCI5VW0Hv04Q27q2xy524Fhj9GWgsUhf6UqeMwJmzX9nQRBsgeRMTkXmmq6
MB3xmnWwp8oUTYK+vSXPvnKu3ctJ+3Me5QHZidCzAOTYbP+ci9iDLFo4qAKSYhbeGmzwfz+NpWes
x14jB6KAoT9W8VX/k3vPUne/bsVkxq7Li1Oy4Sdvao/b2ELwgtUJgh+zfJYXFeIzUXdrsGlLzbQK
AcFc2Ih5h9BY+d7vyY9oYqcCka2VEJbOAEdaC4BYbdDYyIOyxdqTfPO6f4cEzhRle5QGECyuixa8
uuQ3z6slNiTVQX/n9JCYw78qjgllJOcIB08EyoMZqDOI395BGoowsDPtia06EUkG3cf3G3DCAVar
Px2GDg1XxUqNiJfm8pWfaZjEhuyvxL8pBUOdZUQWrmUru8DfVovi0c+SmbHKMJu9WiGCID0IPU9q
QS77xE5jGSCmpJA05ru2ozPb96RxSuTvwvr8JKtY6kkHrDNdDJrgH84+cqTlup47YNX9kB1twZmp
Gr308U+/8QrcehceMXmWmALBK3z0vK/2TA+D7Ts73Rg0nLM9I9VlqyYAQYi8dbmeh3P+pXivz+BS
zq9Wr+3p8joz53ewZM1C/MLmOJhFQC/iNgrSL1w+i/MHEoYwElOym0G7x0+bv87lC/djUxY0GXQL
rfXnN0cAs8Lz8nZs8vPNuSzZVdA/a3X92PQQpN2eAseH1DtdI+IxWAXczB8unxbxas1FdxYa4iHS
txDUWwRagU0SaIwL4Bk6Ceo6obLPM2hdXs4CXhAb/NoL7ww0Ms28J1Q45dLQdpYAPgQtSrpE0yGv
HVQxU6Dfvz3tGkBO2He3DPEfyp8mpGNvZf+TTlL6DlasUc/2xCUuDy8Ibe5ldE5ZNO/bH6CBF+Vf
QJjUF9L/8wTAo0wiwxK3Ev9hq7bbsFCN06bZRFvMUJeFQ1OqeOUBVbhh5RUOZx9DrbqXkxhgjlZT
GU4y2DgRWaHiSuqnsPNJenLvZGKkZTbGh2wRDCiT4JrgKV5TJ/4AP0gyidPuxrBtb5mIl0NM9KN9
CwM1afPgiLB/w79O72GUVSCe0Q7n0ksdDGWxK3VgnBWiFRzp/XzGzaktstQE1D7vPmpuSi7bX/Ri
slTuZOyucvenSRefx5C6MnMnkf7k2gvx1rXmvXAVVyB2hca083omooNoaE+FDTge3jQiyzqVUPKi
mSIDrPoUuaT20w8qW4LYgesDaMQa5Efpps3YL6Cy9PLrFIYu4hvNRpxPu1gXodTeruGT87mC76i+
Bu4P51s564xdrM6Wac1QX3AA6DgCaOZRAnQsGYLlq4UMlhneH4E8DLnYSZiVaePN9PM25bJjIDHs
+Tjrrdi333khC8a3vpFtRMEGz2CXmdtBxpbXRUnl+Jis3XxtFx3OEvkgAUQtZKH5dCckmpAGpvJD
elUVO1uwWWuS7H3SVOlGCZfRjKpvNLnt0JJJXVDVfV9w+xGSyWG711k8sb8Qsi0/aEkKQo4SZwHv
W0wivEg1SCdUe90gHfkrs397FZnRk4EdQ/C9rG1hPI2ZT4t3ZF8po1opayoRcGOu0HqfJ/jFz9fz
kOEmXgZuV1jv9/ex9fp6djAJZ3WfNAt+K/inQlCXrc15kR/CUDo9ZsL2PlGXTP91TP9RDbtab0jQ
FSUml+bJVdbm6DBnrXEXzWgsC0Zuqme5BvgYXnqgwPb8JG3B46anJ95nmd5XtFnzeQ83miSxBfk7
7fIXoOegsXqko096Rzr5YZsU9PjhvTmth7IHKp5+vqp3h5lvIQuodUyyZp6fwC5qjcHOnTRBWlLw
uR6Sn9zUn2y7cXZB272kZNzUAII6mCMNkDNMZOr3NQVKQWqYktRpb9NP9KIJ/qKWBsNn2cBIvbYu
gK0SfmBtRmymwn6gUNdq8t/N5lfma/iuXQFJqOwMuNtMmEkofiHKDoCOXqWyDl5v+I2Wu5JjuMc2
V7FaAgY39QNFHcrq+NcRfOxP/COrB5XrC0Z8PWlnalbzStMchi5j/YiHMcfrjLfCJ6JRC7slbmlq
cXGrd7R7bHcQPt8TUX4hQtnDfWdKHhb85EU9ECMzA+JSPsEXVIIsgwZZWbrlz4v6J3kVOKF8lg2T
pMzCBFNqxR0luqUp8HzB0/p8qHHD9iw4my77LxJs6qVQ7+aoGrWpbgcFNDdBDsNcZDvsLJMQTDsU
mcbNyVQNtGdhOMUrD+3+F+3DSVdHwCov8KZnUbUbkgIP9Qpuqs+6CVjafgfs14+7hdtoNE/Xfcbs
t/zoo+/Tz7vPfLm4+amOZB7oFVG81HhKr/ciOc7rhu0SFCcF1ZxZRmvE4vqs8jWG2NG+UIt7kapN
Vva7S63i8/Pa0X0lceODIjsDmolh/17whwbh06I6AD0d1XHGxOak4iIy8Up2X0IHdHntWTKcKs2P
hlHKI92XuM3QIrD04cU8YRTLDGxzd3rF8Tha83KzdkpjHB5CpvToX8FYn27HpXVPXD4UoCndJG1C
aoFWBzI20hF7C8t0pqQD2hiHUNglaf4D6TW8MCwbWHVfxvLeaRcwOc0rbtIEmlNM0aM0bBiXF60t
8y5qymFFWg6DLJxS+GOt4dpIivD4ts48frc1+ZqZtLxe0KATrEh3OMTIHtjSLs6xNuqU137l5F6e
G5AdyAgzNdMSyWfzEaO50IckZOJo+KuJ9xz6PJM+nRUSBb3mUY32zmFTR/vd5gE5eRZ1LI4A+GTE
QtvzZX2jcFVkuliSb8kr/D/ggv3KQW2Dn/uWNClCunx0ZV5TMU/z9Hj3jDWbOuuDoS8HgFXguqvO
i9zsyuryWmrENu4UC+bUHtisnZW+a7BBysgaCRxeb+6/UhulTp6wIzv0KEMRopXs6ZhZyeNNlmnQ
n+VJpSD6lgqAR0p+bH4Ubm1RifwtWUqkENJTt6DlEpVq303S3YTwp7rRwniqERUn5l4yRHworp7B
P5+u7X+iXZs1S/iyQGlEVSdYRbY8aubMfvNCJZBP+NQUpAjEbO0w6kjex9TINFJReRFoNu6A0/3G
Xk9NMcto8Xc7fqJs2YyB0yrIMqj0F91Jy4y6fu0JUL4Xk9Laqv/v+ap/4Hq2yUJxiuvyhY4JcQmB
BB4sluwjLnyH3HRHTGtxGzB0oC/J3nQUxKHP+ntadbMAmDaYhTg+sPxf5vWntmyQixvz1MPRj4sg
M8zc08H3j9WoUDk5N8HD9izElKPBMpd24d61iYVAY21gVqE2krowXtiuuU5PYO+oY36UXA46eZww
V9Bpn1BhVhM8AGTEOCEAhADdccyL8eXQ5Yb0XpWMg9VTYY70gZbK+IVVpQQBF4D1PL7AIstDHOkg
t//C8u5/i4ZuElsIEs6gP6CwX/Ut7i9ommewV8crL+mxi1lhM0LA6KejtJ3G+kZjANIEzZHuW882
9Es6WPEtTWghsnNvDC+lgJUo7rE2iOvVHGOG1hqw7B16HiOAR+FVaB1JFpKi2a5oV2CXX157Hhjc
WnQkAc/6RulG2cDkVH9gbMghs8TmJS6j2opJZMlIT/OY4inBNif+drZbg+mdRe+mH6+XU87G0qfm
F1H3NXoUTV4xDONtfeLFnTgi5JjX8iIpxUdHL0gqm7GZDQbAknQRL63ZWxM1H2tph+SmfCUWzJBZ
WCRZVnRM7TsTeYGz/0vfG70YB+UYYpPR+XSWm0SuLW7QZKpZ7Gn155clzlISy1O7gOVro0IwvEUS
ok9Szj2e3A8gmqpmCI+4fQj00l4LwnJOO+3SC/OBwtOW1CHZElrSybXLdl3PCZSpDu7aWcvYrykY
ZwiSEo74vlPDWl66rDw38Bpk07iKHU1qI2JbKLLT1DaV1anjRfCIIeyWzUow7VLIOdz9RKAcix/W
Pq/QEb18DHzTDubMlDWPi9vXBdXqwHDXux4rvgKjFVmtbwC6hrNUfiGcp2G01vqVG0kwSQMt5OfP
kdUGUx1YT40n//HWWR+xdQi6aVLdnZBssa2xU5CD9kaCgC8IlzPr41wps83AceK4LhhBeZn/MMqf
zddC6uREYwuuA37VuBL3AEmaogwgx1iVwIcHsWDev6tCBiJUsh4lkuP7MZOWMcxvEBLjHzQjbaQD
ukxEKyF3PEsI6Ey1/vP65n1aLVOyOu8iqWB89ulzcHBeVdNVMByg/eP2bWaJzjiEcf7qP5jTbKrK
OrSplTCECyhdM5H9hLumWqliFU6RYA1EVAGSPz77nfPeQGU/ujUr8gWjbyco3+QG2ksnmLCJEdeT
TaLqVVWMzrJ+jtX6O5CiwvFNj3bXTL3PvulLPBbhQ+E8DEvXujCkNc64HcL2+unnbuorv6wpR6yc
kwcEhJsAjvOkXWUflAZYs+t5V1iUw8WR2jYDjx6TMxpxfm7jbJ4dEuJxKRxf5yZx2fs2FXYKwtNv
RVRb1uNYaMRnEaNeNEgzkKjBea1Hnp0oLwohmBgbND1HWQngjIhFUtGasutO5gqOoquvOWoB7C7J
ZJf1f5gsSwBffs8kjl4NySWVK3w6aXvJOm6h0jWxWJxHnKJervzM0a3XeE8V1CDHveJIM34ifnwq
jjphVSkFXI5Wo6t6JJqySgi9tT3KWaXJE/tA8rTLi8VY7+v9GmbED2xffa2L0m8yAeuRIXDxyrc+
v6q5YymubC0v8tC1Vgwh99UL+OUXn1IldpUqGETWyEc8Z0PAvSb06Vzn0bYQJ1ymvF69HLqLxWAW
DbjFN1xDBhoj1EI+PwYfOEQ6Cvc4zUocG7Ib6O0zEQVmFH0EvQyKfOBWqVulpmYCfZ9YN//3dY6e
zOBuQ1mjgbzDPDiCpf7dDtB3Lcm8KPvVlF60M+ez1xGbMmGRWw3CZTK+qpzrsjbQIXJoAu4XXAU9
uPrBLQ1qldQ0pmcCvjZUyb2c3UaIV27P/iX615YoJVK11Qhvgu8hrUwyCDrriFMwKiKclgV00Bxx
QW60zZ1nwloh9lTxmckYIutJaYmVccmhPwaxsP2oVtwbajVZu9WKQJu8NIP7lqmnslqb9vsrV7Ek
UhSQw331fNiOBBQA/KnzB4q4bcK1oGCGH05VktDhbLPjgLVF+nJJKQTDMvwtMYBoT/W7fIMG/OzB
mMJQT8UR4YVqTl0T9jQr1jeTwqsY2+/mJiYTxH0u0RYhOE9WRKcBU5otiuam+kzVKNpBA7zJr9Pk
q/nfX2nmQUM9UDk8rDql+K8dTFO5KBpv2ZcxiFrET7I6nXGOfhneYYjo6LZ8hnmhoDmlY49u8A/e
UfsCZH5pAWepqBh0/b4bT1QFUOAQSAocvH6vFOnYOVeM2NpY75LE+6JZ1ylFMvqu1IsB8EjhNDsw
hNH9c/BVOh1bKHfDHTdOUlQlKr5i9dIDKxC+wAB0EWPrdsWqgWi8fO7jSG9mVnC+LQAGzGCyGY3y
AfMoH8NLvFJlUPaCj9xhkbceXjbfo2PzMxK7UjR3CDLWrB+ipKbAuzg7WdxS5XyDZ231VfN6FcQI
kgjBfmTU6q8n41FNAf+zmLxKcRFxDJwsDCVAuyqLmiVbMtQBkHv0edqwv2NxfqSPYfKAvuwNuGdu
bo2iFcYngEIo11h4yBi/ktRESbJdfTwExVkxQbab0sdk5EZoelOiwSGI/4T5JGBv4c26KnO87saw
md1PA3d3+zJdPLx3InEnLvAALSr0AjtnbIU4Pik8UMC3RbQfmLH0x5DJlWVd9wAET4owmwCFcvGp
6OYiG7YZLdUDEf1vYTHePC/Q3jweXmuC/E0YKMD315jCGHvKEfrcFwWtlZoqn/9+yb+DMgAncV27
pa7eVyVtcAyVgnGiPBLopCvwbVwV+xSV8NqdXT6OxYhKp7OuHe9/3TqFe/4jptEMc5l/D+v5dGw0
VZ1ATPNNOpRg3Pf3km/UjrPvyyJ9KQNvDSXK8iyTR8jj5/SER9/EtA5HEoavImXApzjRUBIw36QR
sJWohVE9fxtD+CVjlW5mo8zernBiA5yXx/RBe1ABX/j42VlGw0xZxFkR/pJE8YjPSeg1xIgshCYV
qBfKSHhl+TBMxKqRCT4AhgEOX20bwfRU1a2UTkp21V7z8bqNidRmbn5Hmjri6ynqbnTiQaxd+4xM
N/gC/oJ/T2q7RuyhbqqqzKn5G2UfZFwBKe4oPCfMBmt/D5mIlBX341c1WZbw/++IvwXPuWMktpzJ
+8UQygrH2OEbtovX6D3x571HCtg2QSxegrzMgqCvsoz75PfcV+Z6zKSO6OVFl5Ry7VwQ5yZRcvYf
tMtCv4Y3bKNsLxEsKuywlSTRueO8gLUnVoRY3XpQNgVRpSzCr2OIJvd4YMWgeSBX7sjYiIUp1kG5
hB8pr3zReUWdbFvxlD3MLNUDSVYguVnNbiXksDSdXh7yWtXk0MY4OKp9QHMsnLBZzjqwd1J1lrMt
TTc2lKPjoPsJJRg00LOwC0ryhS8TpUU/buQP11QH1kH3el8tDw1SUbg9Bi2onvf8yHTPko3bmxJ+
W5Zf/rQK+rDQMihDblhv+2AUlfzNLCXL7p7XEVyFiqUbWPvc0+OEGu8SYFSfr44tvPur6zc7wJ6Y
qFZpjZsicuAnnDTOvxLM4402ZxWu/anUjdP/xkIPnZFbN75CWwESln+blS2/8eeJDNlxRnSpP3u9
d9VJ+qsSkgHNfhRBvapSBLDAav5VCTIgOketYvB0HXWjYJSnMvYazaMQfbzmzYmrc5c7txgO0Z3B
/O69o4He9OZfrwErF5ipdhuez6McDu40PPaJxyXX0jCw3tJnvEgVKa+39c9xnz+nsPmseiJSvxU3
rvOMoVFf3IhNJ2n8PxLB6tsOIAYDi+SlVd4p5YVk0YFRihqGoXcVc8N28ADT4NHQeIlzYO+9assK
B/bKfw1OH7KOD/XHmlPyKQpJJt/Fym6rrhPmh3zo6BoMGEizRwrFCLfzQ80GAY7iWbx8BOSMEXLF
1ereKuQjh23NId2c1kaz5nGF8Dz72b+dQrS7RrKZXWWgO9CGclWUANOIJFwpSKqtSc3hrqYP++sp
QPBvEs+v5HCXDkXvye/6gaAT+aYKcbZUnTgpsVHobkBxtg5kWH1UcAqRrUfgSgidIW/wNrAxkqHW
27/oerhnVL5D3DhKVjf8G5oBETp5U07D8FZI232rkoi150P/7MAVdzlv+sZMVsSylAAPRJCv5eRW
pfb59rr2mzGo+OQlgUSS39f3hnlJMAoDjARS2hPQ2tQRsrry1gZKF71B0igMNKMN87zZuewd2nmB
uK0OzPJGtYyutb7XCt4ayn2ZKnZX5GXQUGIQa9zKA6piGQ8N0mN8gEGGywBbjW3hwxtW4odHpsqj
JZ6QSIBQci9chplXXAij5XZcv5/MG3zVxm0Ksw8ZQXcRDZMJhcaD2rXv2/JolSDF9b+WHG4lUgk6
eUsNHwHYKft+X72nj12pmjOMG1lCmWMTu0+TSyr4ShKXxlNzX2JMhopiXxfUA3IOCQ0tXVfR+7YH
olq0m+HiUS35m69BYHj3hjIMjxEYx8jzGI3ZjLgA8c15u0I2M+Y76ZKkT86iTnVE/FiVer7jQKX+
wJJKYZFwg/P0/omK9sPXnUXDG3qMWbvLlReetXWNnjFt26Zd/xIgs/nGCcU9f3/yhGmc+3Q4opnP
Ads1X+XXu57BA+VMwXV2IXN+sCNhlueXtXV/qic4v7FYaUoD9j4Y+p+HiI14b7zRBNkKHZQBmP9a
NoaJOuIrxK0FwY5d403MAdLWtyh9/6tchHbbXcBB9BVLAMZMrKyS+eMk4opY74KjExDjJKSY5Aly
4Nwn4fIBja/hR4KiG+CEtnkufbNSgxtCsq3k+Vcm6FrVJzIF30KtFyJFpU6JXKanQYaQl8o8Rbmp
oUUClRnTPl6OBTBS7Jnz+jJdoxOnE66hcQq6UU5LXV3qT7c4rGcRFf31TeKQska+ED+dlJBKIz7P
IZfkTOM34gzBjlbLR+e9yHGg086W53rnoNQpjmGA8lfus96l+W0+bb7l5p2/dMIthjwB9yH4BiOh
9wCMLdrTWR8zXP2MmRL6xAEQTG3DiEnNLhFP/r54oOMkR2j12pAUOZghzWRxiOLxnpJlQDHCi3ro
xlgkOmUcjXlX2QxarDCkT46t4eco/Wk7Jhz8/KGga0cjTzb7Y89ynpxbq15EGHm0BPjeNI1UXjIP
py/sDl2RQ/p6OYjCvsSSwdmoWQmO4ofZSy140MU/SQmPlF5SwZ3hfTZrxZ/8Sl7CQpDPp1u6S50O
ln6w/PsWTMJf6+ePpRxc2Lo3gCCYdaM2FOHGii474Z9IfdzSzVjDZ4IJM07MjbYa5+1v1jEY4u2u
nvtg3gM5k5ffSUCPp4vPxQQYmCfS7kg+Sqa0De/xIoGDhHwvZb0CqTzht7xZkwbznrtLDPSXp9PU
UIFyr+slBji7OhRVpAydH15bZvQXHl7b0dzV+JEoMzb7nTO0IqjKdFRO8xFRsuyBvP7e8fyep/dN
bMi5Z98BZVekdydmwYaCO81/RO3l7vbCzsUrbVXOY3ItHo4tPeuTqqdKLXLyrg/QpJfjDxKN+N9+
QH4tXJTz0XtuOCvDAbtCXVEmSEVuWvKE0tHJvG3DZ24rFf4/r4YS1FfqY8PqV7AuoMt2Vl96/Qni
sUwNwadnJP9BRgGySf2DtG/AU+bqpFd21OaQsj6nR4PZ3dcunQzRmx/qB1/QmRj5ghZNDnieoSqb
xs1BwEEiRH6w+22IjZR3OHhuGRXfmLaw77BjG40zKjggW+4tzXUuzNkl3X8LkLXxyltiN9Jz6JUW
aWc9TdbL/p+fV4weFrAkaAQWVhMpvzpBngE9G0nCMpE1CSgxnCoICiCSGecO1qCzub5Xn9GtXsOP
SSKblh/hjtqsHIRZFyk2RLg7Z0i67lXvinyRGbvmDZV4+fnvNSI+ByUtG4FVrlkeJG0lqhEfX1E3
yAa7QFX8C2k2I4O1vSEt1Faqg1ajfeh6M2NQbSZufvrewyVOgrlQJWfsBVVZ8uOZiuMWrhIzwPjN
RZe+MDWwY9my7P5xwhlEBcctugsqD0yecWTEPO9Pntvgsl6rz8Vo5e8JVPkil0nKTvkzFjTmI9TA
l9aMpABNn6WKhUxMFgvBsVGeGeJEDTkDA+A0gHBQKEeIQ/w3ldK+Lpr9QYuBx9X0iGJIwMhPDzPc
lmCNuxZk1sLIgUw9NUam56GQSJye0s4rUQrBKrazZEUalKEG2QeABewR9vxd0W96efsjncWOZUeq
WmLmjaxuF1b1uhDGgvVVAm/L55chHtOToRYiLkMpPqqPor9+9UTDLr35Q79Al1l1Z4IxiTM8mJ24
MB5E22qtk26X+QN0FgcqtSYXd6/GQvMQhy2hG7etmu4BZWuKP78h9Q/oa7NreFRw40si8PFIySsT
dIUeOeKHyPr4mcNLB1ixGcKY8/V+s9qradGoVLyfVDhCRvSDIsk5N4SVMTw5NTLCj/MJ16NAo57i
T2hvGQ0fJXG/sZ65cwbZJahf0m9Gn9kcJgptcKfwtg7XIVj/2cHPVxilbvvwXmNpbYjin2CmcRXk
z1yj4GMR1EwYcv3qpNim7z+TEXH+b3Q0MM3t2DXbE5IPPAvr/cbiDQHD0pFCI+zp35nJE5GEW9yO
Epk66zw19acZZupo/dexoNhIkj/XsVmc9YZXv3NBthig3pTo2AndEAz1tkp/LLLJVkHlsLlJowXf
YughO77qRmHOBIH0vYnweNZACOnD7+5s2Z4UXlvLz/lCdi/VA6e1n2kT2HEZWPX4A/5Hyu2/BACb
pPkAC+DWj7ashqsGd8ZgSLI67tOZtQt8UclzRZT8pD8oUJpG8uWqBrVbJHSvdDI3d3GElHk+JC1p
opwO1RJweFkzJcUpKwxz6F+6VEEy6DxzzR28E03bISrGoU7FzK3E7AcwcUHM0C1KXHXKieZWSRZM
SXwlXDJwYV3Z0rso7zKBC8GPQGgG6ZB8Y7QalqWfhjqDmucavLdKiDW53IpsJ5kf1hALdR+bnhns
HHyOsMtXf/MS1kIHJT/kKTTWTQbAg4znS0j4qOOcnxsAd8/dd4xj/Q7pN8uRYQ+Ub/sccLLw/G8E
twJKtIduTP3qovflKk8Jf2m3+yEvxoKigQFNWe2/QGzvJTOmCQywDXN36r6PIpYfevye+1FS52c4
LJkmHpmGrQcfsEEWxJxZqtKf3Ve63AIylH76v8B/FGYAe8dA4w9manoWkP5DBHGvSsoDbUwrQeSt
f6vdf3w23p17Xh62Y4HwKSzIXmfCx3rX/Wv8IBaNRv0ssChSZN9Xr8MkDOeSC+vIJuWYEeMagWid
eDKy9s8Mv0GU5KzzRUcSmUmxlCoQosNBJQMToNbMXdAQz1Gd4NY76IJYrZg9N3hGS+dy/C52N5BL
Z0Xog+11hVrdgGu2gYM4ZyJOXqY7NmMWsVz8N1L22EFV+1dBTBLSmWPzCkJlhIR6rKuWqGvru2ni
NZ4QCHKJnWcNLi4f4oAEmgX3Ve9ymdGYB/aOXi4IMVrYvfIIRs+kCjB/jqf0Hij9lKae2I7enf2Y
ZJaNMxLvvZsBslEc6lSmYAKYhW13/b6W/bCX6Q+LinE4eQhtGWdQaKHfWFRkn+/hnjlLaiZLfujt
gx/+Z3TJ4zl281MfnbnLdG2nb7c4HO9sg+kuMy9YogmLydlJbCkGQdqs3RJsznTcpfzbJfNOE9ze
PiwiuAE1xkhO2jDyKJjdSYSHxheMTBNY1aCVHA45QCvFNzvNlV7iz6rqKOVwa/0olXTRDE+LOOgE
bpiRMdwOeFRJpKk3FsaoIGi8iQ4ooDOIBt8liTYivyFloY3RMd07jz1z+ny1FDbDAnEdi5yLf22y
jQeEvbsYwBoD3qp+Irw2Hx7TecigY1rnjXiQm+B1pDuSGDqLRb1tU561wiv7rN2qfhPUNdagLFBa
ND9E7Hu2P/SAY2ALQcHHEem7mKTguh6gBylFuvTN/TjccFzzi43bsT+7ZuGRmm3SlcW3q3mYtO+/
7Fa1OelVnfpON7iyt89Mqu3r+YphwCqm6WTWvq+eQ5U9E2f46MFQxg7Du6sj+zTgzrdAnmeBUUD6
65sw3duzxJioNbi17q1KjfIRTKEdBnpYr7OD6vSVRtPwJ8Lr+Oacj/b421RwZ5ikj+qomyWJ1lXL
iPHrAXnisOh66LMhkAAIP2o3MPZE3b4tUTwuVrK5hlXUaHzxRRcsW3T88MyNYhCflM0PocSnYhOE
aGYmeG++WD2vaXt7Tnn91Za6IJGbkuVd9IfI5hK9Vi1Y92CBJO4DQn6eFQe25G0bpgwTzJT+GxVy
fo3yJQy7evZo6bPPgGs4bJia79t+vvTNHk2B7MhlV3ff2YNcwhgBTmEniOnY3TQ3gXzwpPphaEdB
RBEls9IJfa4JYkQhTOQkqq3FwxOFGameEsxQGIgXa76K4L8hNbxNy+L/zDjq94I2F3FBq9/it7k9
wQDztDWt+mSewGJTZQsTrGOvQbOCQNtnbnVf2Z8w9EUiUrQt2Vp1ewpnmpvI+4ZsUo1jfpHQgTbX
VCkMJAohAC9WPkIxTvrMCTxCxr+Y17It1PsWqXch+0S2y7C4SvKfwx39kZkN9McC6vF5BPuQJ58z
dpFyB9ZrTADBlq1pYG3pFiGLOD3zvYMIVzTD2iHMMudwLUrEUQt2uI06XZA0oEfNCOs+JujCWkxm
AQGN3zNj2nOf9ZS3vG3T08naD3N6sgMIRybZrjfwmU7URM+JW5b2exnAwE3S5InbOzEhgA1PtIHL
e9VA0tRtHoMJxDAOREK3INLKHo7jRl2lxUqGEvEL7qQYKNzfDnHBX+IIjWYPFifi2mpp0NnWmGNJ
GXdBya31RTlq/d8d771XpF25x7ZTleNFMZp/CIch0gGrFqnQ3BvBmS8R5Q4pjpr9GQHDUw8CwszQ
Ia1R1jVsMHWYL0SsbCPQqVEWcwigjl7mzqSfeia3zGW5fwFoQ7sisz5mOjp8rS10+A2QvvCcoPL6
PlCj7EtI/YTxVe6Pg7QgU+E6fc9dmwty64ZNLmtgJs0H8ly/bki2+Qh9IVNaNlMI/wBtEojdQZzJ
UkAa6sZbSzFifx76HLFrEQt82lKQeHzjQRUnNfC3ZrveX+YHe5YfdTJ2WJ62oPKR3NjnIfGpsD8l
j84sHCcmdsLegRL5+F46Nq1bF1K0k8Gn0gOxeMCeC4YMG/9frHMpqy9+dU4BZjZjCrj3tM+qTFKQ
ZXXffW6douRUI59GD6Mhmo4rtwMbeyzggdE74iuPgfBFFSjrvp43kdjarqVXe/XPYY9aGCSB/RbR
3vKaxnPXKo47JYpSJytGLwJ7tSJ+vbC+AfYZQULqV8RxNC+AfdOCuMJnBZZ/ebOfRsKmnqtGgoP9
tiOAnfIwzExwYvbMcNNP33wQ2vBqu/cI2aRHodDv+n61z3xIKg3h/0etiCBP8puZgKBGAYt6s4Ep
cPYjmFg/HrO7t03sWA8x1W32S9IPxpAvdCwwScyagMGqZlwV6W4dtxaJM5kg9GtM9GtHU2RLT/UY
eGsUynMkJ9VGGQq7szRZHUh6eHoDkI+LSS0QtGaTOujeJ6AJ9aHmtzyRhRmphDIFVV9HO3tCixtI
ijrJWTUjS2ES4+7PNj9l8Pqc5mMrKhthuOMxmQtftluqMmlYRNz0o2p8tp5Bb2QmZ1nk3zhWLbQP
+Z9aKbm8bknBMX5m3UY6zdnt+pMoOtF4T6NlBZs84GtIcZX6To/hTn1KV4KGYenUCEFBvB+ewhvb
t5bTtSQunZV7+9hu2OqH7Co6wK+xQrS85WKrvYvKMGqciTtPO8fWZ9UlyXXHwF+tKiz92ktxIrWm
x0EZLWn0LF4GIkjiNkcSY+tM7r/Lg6Ex1yYUM9ihfjKhIQnsCdclJUzaFgS1qbDPqA1i/I8TD/Zp
SKUU19ksbMwZJWAUDtcd41ylhDLTBIX8WQnHT0VcSOmAzMAc8M9s9cuUeyalgBQ4y5DYX9oLyAbS
EK/g/KeAbNGgsDi8SEeiIQyULAr8QjyiZI7gBbhQUcdf4F+Vtk4M9LKaa3T8WvV83dGnO15gP9Ny
aEQDAvxjAqMYIyhlx58Fupqejuj1jczcptQmih6hpniWCVwkAVAmeyJRiAEzRbsWPqJZtxddW4Bm
4T9Swdlw+YGTwfB4llw7+LKsTYM7mE00f19MtQwLeWxF9YR5YuF82ZCqj/mwSkWxsLGH08V/liOM
zv3WhsYSg+nocnK0eQ8M4/QtAR2e7E0Zz2kLO9dbVr7iyFcb3W3COfyEvkDLl/oI/hWFDBccpU1t
n2jlStEGsGgUFMpIED7KvEbjkB9nxuFfER8wNQiWrBQ5/vjY4CKWnEjUQm33lI1AxdI3q0F+JEyt
kFF8EBJD8J7AzK9Cq4xDajh0TTGmUC1bI+yE2i8Y0xMATGjblRdAR+fH1ln8G0RlC9MQBZZIL3RO
WbmZ6rEmFuNWaj0llfg9Aw3mfo9DLpqpOWQij5z4xabagsPHp/oifbjBnc9pJN97ePSWznyoxTJe
A71Gg46HBu+n4CzlzBQSIWOXp+IoxXrUKYztjkQu47lsmieIAntzEytxKI5NGa+UHBr8jPBahf8B
dS1Raxv5w/1HcTDIUnS638ApWSR8Kmfe5FS/JL6WCYkSMvdifhn0/KL+GmYZah8NGtfZi5u6l5oV
N/O4Nt55BV234dOdMTuSGeH2LuJ3vHuDP5FMbUHTRABnVvg3W1OHNG3VVqHS/ujXcBb90Topqmoj
459eCpN+mlWPinoKhCj0lPdqCG5INUmRozMzb79lgwNbAv4BmMneB8/e8NhugRwIfKtuOBGiorB2
Lh9xshLezCkfx/qCItw9enEtofoAgItlXTRWKcJ4LjP8wWSou9hFyLIRBvY1z1xW3nF/V6BQhzOD
1Bnemfw7ibvELNZBpOdX5+VH6bomPtxLaEDVmFvpsAS0j9iLDAZ0Nog5+sBKUFq9IEzlnkooGdBo
FDvzw8piv82amqf8Jw3Sq0NdXzwJekZCMMlJ5FPeI7Oaowhp/TkdADQOxFYfnfdHQ27X9goEJN7s
Yhz0Ql8xRA1AK3m0bM2M+pC1Q1zoU+SCFPBWDHq4NbnX3QZ0xBfJmEA/jXqIrDWfbdZsRiqJrQ7T
SCggGwQIaoH5glAFp0rPc/q6NVE3f4Rm8G8To9peUDNGlhotaT0vMTSd9fLPnq8ZQKNm5Am4se7s
9QH916+RwBOTiyv6JwwXlO0drhb552CZ8PBWvsH/SALRj0d2e3Flq2lwA7RcNww1l+wCIok0Cqmj
+WOFUHNKIapNX9WsxRLeqVSL1QAZMhiZZay7q9VFciv/mwSo/biYcyW5Dff3PwrNF0TmJpfn0rtN
N4rmhyOT2FmcuHL5ysHaoNTakZUDUNBMetgotKjL2RwB7X3xviNFnmccGd+w3CwU1/ggs9RMj89T
pQw4rFGge1Jh0ZuoWrh76fEoq2LnwPmbNM+n9ehDhabPh0FzDSPpJRNWpgEYKDOG2CzTXCmPmaCk
Zrg3ecvBykiTjp19yeEYi0dB9r0VXXRB4zPhun8qZwJW38dkYWoZPMcpVY7sR3DIZpu54QWlfKs9
3aAkvTDkMpL/4fYWqnemR7syOyrjVXPgUKAXGDP/iFp6oF9nrQlKCxRgxsl2GFONyRHs/BEXoQzu
C+1g1DNnhbzDsf62jGJm2aQeoqITcNJOKFWx9cW7i+Fn0btZdrlSNcMAPXgFXtcbLqu426XE/78f
cecDWaHx/xJr/GQu2tSFrFTWzxRQy5GM9KQQZNgqg68jVD4jg8eEKgVa/VlMjqeUDttXFLuPzafu
YYG+W/wEJbNovkgBEW4/O5kATJwUp4zZprg/jGBpBSTvwtMfWLt78gt8y7muXNcJMADsEzMTuiE2
goXplo1O6fw1f2hhwtoivRSgUFaHarEmxG/f306/CCZkrDn3x21vYkRHN3FvGpTUQZjJp7wgMHtI
z+od7fHxRdZsuD1r0JWZ78rc2qppc01Kgwy/k/4BoN14XL6uWPumDJ/jT4zqvo9KVHUxlEPFJ3cD
6wT9CXClpJtx5cbdRb1RS/RcSfJOo87R7EuAFrp61YtTDpz7R8sqs6KROoHb50HezdwamF/wNMui
xKEIVADwyDjIvXCp3evIhMv5jw7I01rDo9l3xvhqqOOjzW0p76ALdeBE3Pp9cVKL0ee0ymBANCmv
x+hh7eHwc6P6jppnTuFWUA2qfHsEyQtul5civXdE089DtjOJ9vGuRLXuRCCDrg9V6lxu9D3nFzlH
F9mCCCN8+agAhFzTE2imrNlMFg0xJVUHZWoREM9Gr2T973twyjIpeHc3FeEEuELcrpsj5WjO+9Yp
uaMmlI2FiIAO5uEc+XkyCF1/RmG4uORFSrcGozbcWAUB2Ck3+ZL7Bs0cpaODDe9oQfnJl747NaZZ
LgtzrjuvkazO+QkPVoUI4z84fNG/srxmdHPtDGViyfjE8YVZPknPYoLEz4jMRr5irAbX0Fpuiyhk
TqbunvEKPkSWZwV+bDQWRDEJ6nGcYGO43ystfDsPpctPf2ig1FuWB+9DYl87pPvrK9p3E20pV8y0
BbzWNDM3xwosazvRqEyvRIjvAcdbgr81sIEjR5d7ToBhFOzX1XEE71kzaotrJdPGIKqyamReW6BD
DBohCri+ivuiHlnhLXrr4f0d8HwsvHeE1Cx1h0MhWn/h2YKNTcLzvb4gK/vePHXKSS9eWdFX+9/F
PxB3/YCZDZfom9NnSq+Ko+CqWmsyX//xf51vpmXxL8zJPSWbZ05AvacIxzcXCEOyeyG6M7GLQT1B
jiX4JtVNY47gq5ebHA6EkaIOBciUKGFdr8gAGv7/AUHAOtYk9/5skdf6b3rjf+clGUD7POdCOsh7
L+WKD3r04l+H21NlfXu+NJPtpie2QeA2cdhr9uWHVXjb6KeAobyAdBWtcIQPJfNEv7HIY+pblvaL
rqc0zRHAU6xu/vmIotzhPlvHdkmo45Owk84btLI+NXpG1LPQTegLowkxPAH0k6wjVb2YuOBLZq/M
VLDL8ZgjTt7Zj2RRq2wkoo8jWeEer4NH3C7p4/hhECr+vz8mNsdAVEMtgklW9CCCeqs9o1vT1uEW
6e/wJmu+j4V7cuXaIALZJGb8OtMXv7ht7NO4feS6k8hwW+XKU/SMoFoqkY2vSTcdyZJcN1IS5cWk
XzHwTH+e9xCCyZnfEFD7nANXA2hFnzYQXz2yKXb8BerrKTyB1mmWa7vnAV8nxMMnTR/I4IRdYBLw
a+qPexytL3+sQJ24qVBT1j9FVWsp+zTZ6V5BuaeUgPhSPsID1yMbHU1Br5ACVPvG/IG6oUoexyNj
8cepHJcFwf/qqlVp5ygODBQXC72woQJnHm4bVM8mKkQYvVVbytj0ayQsFr7303EIBEHBIuxhi49t
qAnidhh+eKaPaVZDqY2Sd8EwWKUu3eMrHzdC2+1t9D+7zvKVF6T2qUqboqaojCNSpjrDwwONK2eQ
/WmgwQ/j1JVcEkaGdzruAjHiPQ3X4fV0pvSBzvsK0q3Hrl3KXQ7swmJFm6BhxEfdczLn6HQ5UDPJ
T03rafF4cvTcpA4IlBiu+JAF7on8VYFX6XJa7bJVvD+7mc0QqbAANwxceJ0R8/pum4brT3EqLDob
wv0F2vABN9CkaNV8nNbnZAKGqjxxLVTXm5EoUs+EYhfzGy3VR9dXXAFleu+vTVIm0GMxcEydAADZ
3XYYDEyeIUfdLGKZsHzSz16chNNkBE0swTFkBKQC/2XZbJfwZvW+ujGrGJnjIfnW+vA9UPNfO90/
jIg+RCYuPKmOI1Xu0VV6E7KGDN+WSsAFLOcx1+klo//l3+WJZia985fmuEXzEw5zsfjzo21l4fBc
cse7BiBn5emCWbH0HIrOdzft5U6i8BttR2NCpltY1Z5zuTc+QsTHjPX10wSmYGCZyvHORHF0ABdo
TT77pCFg3JdBkBifxsOUjN/E2Q83KZdFTQ6iTh2wfehgrnRMet5VVO1m9+NNHKDk50txG+Dl4WQi
MkDhi0py+vLx/SCAKalGCaIQV50EQBI4/vKYI5Q41h2MjHeBp5pSVmOwrR7ZKvFXkzHpgYXmoafT
r7rp8kTP4PQaYLeakgE/GFxEmmplXTvm4yxi15NZbpIOj1Inukxsq5g9/ZU/NvAv0Ow+OiQrwyHk
o+K2iPberJltVIEyDfGHZKiVLVygESqZgnUxsD5sfJw6CYy2V1snXm0+xZ+JBdzDxePEF4lbRFYy
Ia5kFxn7cYQgJdFN4/Z7VUPwAlK6qFabylpoxPVmeerhukkFBO3s9PuqKRG5yUzpYXx35//b4/mO
GKh3zObnjfYxP3/mKxMzpBXihInTNFmwprEkuAtCgSJG3vj91Gw8YwhF8KF53dd4+Dwg6IPP08p+
cxZn+ABAHJ2vkSql+kh7f9+5JhKTfROIfoGhfhUYIUWXP1St5z0R6fG5LMdQgVoe8rI0DBdlmmYH
TzQi7BIlIKtdjEcg/u5yismcTAAV00imiakK3ppF/B5kaAjYWU1gMJTMZ3RRaknzfH25A+R9EKrj
ZjIJKswopxg0johjy74CKuB/E/+6C0roWeJmzjB4cgoTU5OQiOwulNi3HRkJBc4cbgFjnmltjHHu
b4DCWJQNBlGPC+OuN4rDJdrR44YDRs/lrSL3Z9OB81wWQUQ/tnW5pJ9vjMEYKolHng5ZkaaSAi32
SR3HkC2S4L+RA0PhbhNMko19AzWp3qXzrJW/YTBPDwybIsNRUCeXG6LL9f+YGw3/sLlB6uEWZl9r
e6BJgR9S3JyWHbegln4OZD/M26vcA2mWLGrUX/sYYZI+Vs6kakt6i1+w4FbXJ8RXnNPv+JcG2jNb
EZIW/OvjDVnqUa+VaWki36PUOkwWaczQQqBcMPosZB9UFVjTR1fLpSCSTCnnbaWyBY//x2ZYT7Ce
bhJeD/cp1SW+Unfbc5tsDnkJRkkNrvaZtldBQz6dB5+IoPDkVye74oSLcFDNvJ8qSaJjQw8SVkuf
7zdMz6XZ+sLjY1UgW0IIZdAO9aOItaBl5h/0gx1YpCNX4eyz8vREi6D3tSNRXgu/420kdvBwdy/O
ENTKd1ztLQsNpjDNzX1Uk+jXC08X0neIwgwScdyv0m2FiIVJ/V/UV1XEc/vCo32HFWNFGauHRkfY
Un5HiexT7D22rt9kIzgjPeLji66mYdEuctYTHdUAKzTBueUli/Kp1PJf6wcBeqAsl5bEbFnEIn4d
XE1lyM8OsjvCGnqDZKQX46O29WkNejRFpQO1ymWjt66UMsWdKBj1X08npHXCqx7CxSF5CVmSAH9V
K5EhKbz8Zn/pGR0fwNZ/lJfgPCudb7glkz2kMwaMNkYmJa7d/vFEntNvUidmnSTgk7Mc5TPJ3pdh
GtEmtc6i9SiYpzMgXlgjosLbjSF3n6dPxOKw+/gWcSPITNKJ+IdX7WeY2CgjDKNW6Tdgo5QlAZkz
zHrhmLyiHNB6WoZrfhwhn8MqYySoAQjlOl5//18JMSI8xpIyllXWU4yeSOGMj7gb4cpGfsmCDCoZ
PFVpcF52frhnxnL58whRWEtyTzNAg4lrZpt1ug1QbYb/YuILoLkS2hixTsR3anzMzP1eUoWYZViq
5vVYrlr2AMaNhZMis7kCwuiC5gKRY+YJmjybFEGKo5ifQSomoldWCrVE14DHJwHIr6Jw071wUQz8
PJBVJ45t2bOxcRYM3i7CppXlaei5WVQbV7J3t1MB3f6ZE7HpiHfGak4M6YUwMDMI/b2K9W0SZUEb
tNJe86BZ/7ppACpJ3ValedEalP+g0N2tnBY/HnXumzAR9gXwyNY38QLL/uEEIQl6dvtW+VF4SHZ3
iNg73gr6jxSEchHqU2yZlFVxRfij7IR6Hd1gQit4qqv8KiI2VbOAsXbX3pfeR/K17nt9eqYnCM5y
K8KEedc3ezxXQgCW52cd6GUrw7Ak59LsqS5y6JH1SYNAHApiimtaX5eRN2yVvDNtbjGjnW7khKzn
/hAUogHkMUegp2RtTeoQ+cLiYASkxyVYRq1CJf8rHFrfAJ4WYyxjV9xh1ZY7Y9dyZaZJ6ROOiHGj
sIC8W5+rXhveayknE7PDGg8pXkRLoQYMif3HqKsnLx/ftTjCFgexPJpMi/Qvm2IAsS5EyHTJGC+y
HUOf/JozGudeLsP8pNd61EEi1Y4qB/iAGZUnZIJoB0TPwCxMB+VJttb/bP9Y/e8cdCf6bVnORsp3
G6UvTH2Yc52R+i11nrN+Wa5nqpwQPUZXvvM6O7ejztUrMTucpn1RyLYOmFZE4mcgN0OMy7G4j3tG
LLHefGg4osEMp41RgypGyml06yg+apPpEdEKh5TeLxZ6mYqDT5vC9NtH7v1XmCE6xZwxxOEYFEKv
brvXXkMUE+a05Ml5RpUWdLDpX5eKhRaDr9SiRl1GkRwzJnLq2zaNasskTME2bxr9DjUxid8m4cKq
w4t9akH2UN6L81oLOYGQTCBKFWAFdpDDgLAfmm3+LNWUbiuv5s5mYBkBYIn6GbF/mi+uGz2+aiqu
2qi8GnzkIQnFBsSF0w4PVj3kr0zeZcFNIsCjM5MLE9I9EqFXubMAChAQK2niX3rZYvaSjpDsKm67
FHaGwPhZ/QCKC3K/91cfvgtzoXW+SmkjP/0JWdEOmoU6TYOQKRyr9GFfGEgasx1GRnxKZqMFqigP
XcuxFtx+wgsdytO4kolWbV0mrAr9djNfzkF/m4Y/Zn/Q/fTJuBiev+N9ST+E9UarDz170Rxf8xhB
klGIDGPQrEHN86VQmqtzH8lcfzrMEEV4fx6j5286Tgb0MwRvGSrYwN12RVldbab9qv3AsMzBo/FJ
3v1hp4tvHIXWcS5e92ze7ogHteKIt54KIRGMmJnLKfe6bouI1aV9ZRBe+yqWT3Kodjv6ckOnET2r
zqRu+T9iy0QE0cUzMAo3CrWoSJD0WuP4/yMLXBqnkX/fQQC+O1Umemuw9e8GB1eUImbL+m1iWnBl
AIOP4Z9JDCUTXbzvU/NANveNY77Vz0ajhX6ImsuhegzpwNBilyIs6zZY0NgdNgCiExaaeTrQmvqh
AcfyBHZ8HmSi9d35k97SAGvEHC4lH93mzx1mrueyD5l6F2rXo0Li5tv4pEQa2R6OnOKVG3Tu6Ukz
UagCG7Ljf9r9uzWcW+2SrbLecRE/wNkgEItkiJBwtM5p7w9HFh6mBLMPdyKA2bfPbvV2qlauSQ/A
i0qt+sf246RnEo1fiW5d86RQj1XxXQ1BgkuVbLBQBJHFtNp57NTeogB0ECb8/PZZOHmbm97aDx5U
bt7j4S+qr6nTLIs3+6RrZMWQPJmq3Rq9k2xUXTno7Pl+Aj+MPG1plrTDE84Lu4IOR5QZaZeDnabj
MbjwWRrTi3Nkia//9Lk0xEZ7WMvV5CTDZAAj8QAuzUMcA4aTkK1trYT1WZNze71vFZUpaI0kzexV
a2DQtfkIlNaq07IoMciExlgDrtR0PCfLq6znx6EMd+67rkniUb/oJVlMik89afyEFwzO+AgIKGwi
kk1JQuKzZc8RapgvZgTf2zXht0tOEW39saGoL1FAQTlKwmxCEUWoiQ9/AJVw0Jox3YoKwU0hUMyg
806yfCSrTC36t7ZvqAqzQSkcdf6DxvK0DhkiQVtUA0TpQpOAP6sexz8zuUweX+uO5v2RhrWSFN7s
EROK7xhy53JqswXrQswIMHS0T9rmc5L2DL6nnf3cTXv4JxiaEUOHrWXe392lYltz++8kpPZX7B3C
HHu7vOTwTs6ZLx0GrpeGw0YqdYLXndLpgQEC4kfk0QpcUfvYh7CoeaP/6qvPPvb6UrXooVgpsn58
X6mo4ljTIs7BRxI0b16pfGZZwbu9tEP0kLhti6u04ReqntUU2y8FJ8mb+JRoX0jTy/D5+rjXLioP
IfaDQ37pXLVuZwEpx2sqqfWslNuR78hIOjvDBKUBh4pNh9SOZoSHjFp7p+ozxkwo1Jh/bWeQwv6Q
wRprHeHlv+BczoSPOejK7BCq6s9WXwciQ8IVboepSQIJa/hOLyVaKHplPbrWEFJaOovT5za3T6/O
WbgpH1HtaOcZae6xAB9wHUgc/IHNmW4l6vCfa2eWDy93vBIOj/umyv+uTpDCR1bjGLAw0goM1S6R
wszO5/6oOpGmRM/BLUeq/FesRy6A1v1Z3h6jJDsDCyG9zUnsYL9YVCWAX+vpENYOcvo3hecM5rUK
lgEF5KXAOElTOJCfLsKCZs9qLB8sKi52FdyF0SsfpoVU7X0HG4NQXfcW91NLBaaJ68obgu/z3TFC
pDNG97JVjE04P22OFxLyc6soRVqCHynf9rto3XKu4oa5poKF/VnZH0zPkzyKS4bWRM2HTofsV0Zj
XJR2ZfaiNVzNFaPVmkehVT1WAZDgJS5kwlkwNZpku8NbzWcBGwExB0y1XEmL4YZfvBHDGIQMNbNU
6/djj7LMsXADl3lgZj7tRJuoVEnCIkSnr+eh+hNUBNk/CK5uJ/OU3nztGLhOD/zBMdoiXbEQ12h8
jn6RJKBuI4Q4oGYV/WSDxAMBlDGt5bZd7Sz0KR7cKHhOxuVWMp0gzW0Tq45IAMy7fJaqF65CuE2u
D8ZZIDo96Pj11VZvRLoV4C5zNbABSplnVj06MsvcZeTtd4AYsfV0xnpVEh8TugMwXaC4iK1KnxDu
ecKcYgDaMQ28+GYQ3KaDe5A592TNKjMgLDQL/nKTt4A4Jjwb827JSCLgTVbIq7h4Z4KRrZuVd3AA
1TdVfmgrYak0h5oLVNmqB0Dah78J030sSuJrp8dhWcGVAHMjKJ4Y3z+oZf8rM0xbRJvOGNDVDdDj
/ncCOrP+fYAanjZ3KivnygWzFra+sOrnULSyPcYXNjZgsjFuYn1fARYrbC+MAwSbCBi87+5JGFtd
LnE4heGkl46+boX8C3NfPgfjU+TIOYxbGhQxW+WsQeqZimlrDXDOw6kTYdoV4NxUu4zSAx2awO6a
yXtUBaSo9LtNjs62HQ75ZJMQ/ZfMP+h+NDzH4aJ5Fx5znqd7sJ0O3Cnz6DbEoPWrW11lOTUh1vB/
tntHXcXQArImxIz2QTUVwayeaWO0+gjLkc9y8nIRRI2cw7UkVx0xfjurRu75aHWH15GxzXPjauGr
BKWfgjJ8Bn8/VMbU/TjaBIyTpK2VVDAMg02PbbkQn9F1OFiRFZwElhdVyy87rYbCJFumxNLV7fMy
6eqa2rC8BeGAv8QzFtZY05alN/YaBwisD6te7kl4cmHRjs/fMmHzqbmBVNiII2k3ZngQzHaONuUj
7ShEfUi26oXI1Ep8KO20s5XV8+apVBYJWISDU+MoAPlwuraElowDcZBOV5BlhN7v4TGh7YjcJix8
oj3OIZZIzZPsxJrWpnCBk646IYy1xtYswOpfn9OxRE+NRUVrA7lVEzu4rKOc2nyQHDJ6GU7DMJxU
BeJCNHrKKyCYLM30L9JZnFNZrZ60ScilQOxwOmVBG7qVYpSWY92UkqHDpkr341CBgJ4rfN7TAZVq
Dr3F0rRyChilFH5mdUVZmeH0UCpggnqseuHbVc9wPlW3WsysS4egaPi+Ps5H71zmntTus43XBqR6
6N0CDak2VIew80U99nJFQl1OE+E9Y+3ESNwTxM7v0WLELEeOmSVnbSV8rrLec9nvLQbL3GR+HHfV
77Haz+Af8Oml2bX3Pnlah8TYdjOAgCeT3d9/N072HwulUGu3WRQgmeFEq807HZz0ej59hp8e8i7D
KIGJdMLp5pxR0lR3dlp0sacaqF871tp2d2okDLt+zsfYmWrYMm9He5tvojxObx0fkbhGaiujPuqI
MfRHajSO+DeteEROZfeiYjUoLa3dCLS/YRdBvAmNPTlVqqIzJRZiG9mEt6vHYgZNuaZzsJtoa8Zm
ITwp/DCRmowSPKGc+ujzMjgFJTdpvDVNDi6+A59aiS0twAm8WvxlQ0h+fVE8vjMK+2UhiE6/eIQC
CjzVUhJj28CkBpzC9yPSMIyRoZtJOoCnoErtDuKFHumOen+mIfVAsFS1nZegyrXRA8+RbFCvYx5t
GErsiLEJIC98leB7Ar4l2MTFB3x+qJL97CWCj2OyrVZVFCNuNeqGoM7AkU2Kh0aipwKUflZ8NEMC
x7v8QA9OHvAgM6tw8ZMzti/k2RSszjJjVXYEgtrkLPBPEnJl9zJTdY6NWi8qi2uFKP/idarp3QY4
SVd2Q5zgGW5p6YKNchOWDYwjcyIp/+h0gK61JJfA501gC9kYRGQ6Ui9dVbSLxnWRYWxKjCkiewaZ
+RQn0YZQsEUWA+ZeNDthtAqP3Nv8C+PE+rhUVGDQyXRHxh0NGo1cfVI31xjjhK3g11ZLw+IVw7V3
CSHym7qudO5IeViAk19RNWrICxTa/V/4meGsF5DHzfZGiz02DYZUMFA3UmPqZfLKBum3nZ6B9OJh
chhZZC2MMU8h1ZtWkLWjDwH1hGv/RROtHCsqLTPZ69qgHDQHbcjsgJoOScL9++rP0EEYEL2e+Ybu
lOxYKYlOA+mqW9aAhPAsnfSzSZZzFK4/TQIKm8IQ+SO3gFoVDkYN1nXllfTHLpKgUiKyoCACsswD
iBzysUhZcoLN9ylpJxdiCr0dapq6O/A3d/wEXcLa97HAcGYVXm5hWuGY7AAPcezmlZiutnDh83OD
xbFcwbJGIDzLZDqA73oc6M8ixw0IhFTEcL+pPe049vaVzuFyqr8hWqzdfsYBgQHvu/tzm3hotCDo
eXRTNBxUon/Ky2gbb0nBI8gMp2ODb90bqxqt9reZB7EAFA2lMtN6mXIVCP/kzzFvDj70BycBozg6
sUUf6TR5xCJNSJUAQz7qTUpMD4QoMsKXiUCXDGHGM0kcT6KZKXPLjLD+ok5ZsS9nU9EWU5ndl6hv
E8ecuocaf04Ipp18On68gl0tBn+OZe3lrnqCZvc9xAyWCOAYsetwvrwqibXR9KHo1tQ04Y4iVaV5
ngwzS6CkE6PjX84bo1GJr8xarFUrNfhAH9XRB3/BIZ+fYzFNrocplODotg/g7LnZ8ae6ZfE+0BMv
b+LRI0Akr2V+griaE0Mx5AhQX99S4zJa+j6n5sndUtWQeLmpP6Pn0xzZHxv0Cv/agmVAFe+YibUo
tIu5/Eo+1yAvsrvDg7SFye7/DKf0XmivEWOD0pfUd7iUj9A3f5/8RWqSS3kPh2TMk8yEmQGH69oq
6ISOi/NRKQCGQUbQcKvqitslKqx/qL1rxtOOTT0XfRbNK5Ka7lQgvRDZWOhBcyh3ubG94g6MPMOv
avaFcqImIidc6VlwvJclF+ujFFXc9EIoh49PqWqjR+Z/fPSR+//LG4rVGQxq+Dd/4IIePk9YPyvb
vCnWahJsPlFnNs9yVVZ6tfGstM6hLGAME8fDR2gvN587PTwrCedGXAtbXyFSz8PZ2atJzh/UmO2Y
7e0thVgtc0F42r8qp73Ccm/PBSp+fgOM2jihXBFjR3HyHuyrbTJ2rqaoy5+O01DuL0VfsgrkvccY
WIRjh7/ZZ0NCQsmRz1+pEUVbQTzZeHBUIRXFOX+KTlmJc0t8AWWKFF9wGkrPOhBpSi0ztkRBUv0X
kMXgePwtlMGZf0aFgToC0cBITnmei9QNe7+VqTJwqCnT52fe1HejUdBlkNObOUJ3jaQZ3s8VN+x6
QUfXbP2pU/GHanJnSXFzE6g5o2CqHsQhx5PKaYqOFbf8XL9QJvB7R9pPZjYEdex+GsRV64e7HLVU
SwQwFZRpe+vZ5kLTNCKiu7RTOqFG++KRviBCF1QjWlFzZUNUpciunNDzm9coY1QilulaOWklzuTq
8/7pVokXI67dbYs5yQOqzJN7tSgZtfzj4BLzFfTeMWlGWktNLWUjro2NFa9nKUqLUOjC/4UY9dwu
R1DenAInRy9aAi2Ke1HrfKxn8u8PsEx51DEBN8m2ILCFd54dJtKwUlzfyE4R5EerT3h3P+H7nnL5
+TOg7e+/RQNe0CpF8/kSuxSKYE7L7NqgL/WUkCBxEdhpHQKi0Mm8xgkr7q8WkJhoq9GbR754Db3G
Cp1qMbniE+FVbmXpJ6r3mYxbteirktXwQYq023zjwcDLA7Bke1MT2ymVHMxIOvUz9pCdvOsD7TfV
EZK81GI5r+4Z5KGetuOaAWzsod+pj53sKStN9XET+OXakcW0KcuPpnlNyQuPj4t1yK/3CL4pb1fd
mLrHmKnMM9gvx3kFnZuXNL66yjxN9dG0NDs+x3VQ5imz6vgbW+FWecXZYyNr9/dalprldUimZkC/
1epN1AQmRZPcRPksMflflBOc4YdIsWzn4xnYmBJl2gvQ6BXFMWy8fc/g+jk6BqQiBmB1fQHC3Y6c
zvUQ1tTVc08Z1MPGtwc8rfJoEm84qRRvrHvYnYYcnY3hoGGP1iA/DxBZuMLyMOktqxEo5GizWwU2
XcNjGoGBlSSMyz4jqWmFZQ4hcr49Zwg14ksUheJOXV2oRB2x2l83KxOMRH4e+oZhhcq3q2IlObXy
wS5RJRni7bZG3rZFGrjwRAAtuJnPm+urbdNRmbw1L1+iGYBVfJKoTWitloqttltUpdWhFG9Sh67E
8Ru3X2stiDXoSkmakMhGCy7IcTa/RD30+n0kvskvoadQ4HjZM5Umt58lzP98dA4VN4hEokThtF2B
5TovW4PPRLIYfntThRmvEvww1+Sl0WNE7G34w8WucpBvfXqytkz/9HBSh0QIInP/y2NuNGY+i40W
snM9KelkMS1CJsCA+gCihQ/aS7r88VR7ONSkfxKYWJ2rRAwtoO2USuREAk6e1rVOT2mYfu+ifO5l
ntRZ+NmqMbHd1DXLhF2X3xvsFGzI1nS3iqnqas8FoVUGK3n6+16HPmVy3D1gAtw7hD78GHkunLDK
2yUtmeBjtOXymceoE/9w97hN2OfSu5r3cq1Afp5P+yNfx1z4bjhe3P+k2Y5OlwUga5qTA23ihXjd
amqTy+jyi/BOtzrWhSgK6YlwKsoq0aIlNAA43jl3DdK8C94U9RmjWB+0Em4CCZsvGRoZEqlLHkld
icwpN58iwQ+IbVYjquoTRyTS7/yMbsOxk6mDZWcZmufRP/eDEsuv4ULfxAbm50oqd9sPC9lOv+Y2
DTrt8gx89WXBVZlZt4ZvQS+f8cYJi4vglrrU3Nfz6VQ/lhHWonK3dcamA7PfA7ZrlVKfbgiH4CJG
JpoBqrVIhuoObKJZ+/jZPnM5IjRDdHIMoKBvvAnt66s2GtJ5dfcSD4GGN3dh3fnpcYvnLpWUCLYg
buwc0w6M4Opek9IMmAbkgF0rzCCJe4D3iMaiE+vrlHNT0Pmr5advkDi9FdxCskwze6IjR8jtTZjD
FXvSelD6bPm+N73LbtqdKqR+fkFn9BdcqOHiI1UsoCmuLFXunFzkmHHjdmnkJ+bep4/nGy/T89wc
p5YEvQ10y3SV0WYhHLcC1vfknrh0/kbtysvqHFIn38mGbv3rcLELErhWMTt+KWw+3b5rKwCmC95v
RiXd69eMZaBfOrXbmRa5npdxkyFh0cR8YwxLVCDa2Pr3PA5ukoDyZ+lHnbZ3Ot6dQ3UfiSjh8xmn
+G7+U4Y03jz+jjbBS9qBoJkdGR64UQho+cjRs2yiJV8HTDwrbz8YJLyU9xnx3x//xqMROLjCmt22
f/d8kTVeJpFRxJPasxmuHTVqf0Pc24aq8O0JROvkbF8nzDF6b1y5JdFxqnZSzSS/ZaY1f7YMIqwp
YBDrdfcDGEVKJaMOTR5OFdP6j7+nZ+iTRylLNPWHeIJYd4f74ZvhzCDS/3dJmNQYngUlhhQbx3gr
2rqjsPtNRnrI5Tgl/L4+nmkkQM0gQGu5XsRHb6HH6xMRm3EWVFA8AciXq4QIUPTSIfUWNPOj1xz6
04K4fio63X6HLVXQGOq7Zmxy/njkHuERP8uZswHUOFIefHzZmfX+nIWpOuoXL4WuR70n83U+BYHH
5G3RF0JUoT8y1Vzbgkm4y6hIFc0CPFJbPWxNbjxi+C6NEGLSsbKeJ/cRSVyo6ZgAYGS2NnI0TSQB
HNujZid7vjdUQJ1Lv6aPxy6vb0iPVg2IXa3994ZgJT+gLCYFGK+/8aC6CEX1eXdoc/wVF3JqHKkb
LP2JGyigk2iXdOu4C8ujwj1A0pMgZyaPL1mN4UkPSU5FVsP5uMhj8AaCYmDAu8Ck+5ybP91BjQRO
ev+ni4TpmInz+yROc1CvV9k0UD2gjFQ2lxTYLFABo/wxo7I5aEz3YksPjR5/dp7gVRpSeqbrEyCD
0LnxIPvn0lEfbDtUeTYpJgaaBz4jiWvmRFhae9ARjnbar5R1S6ffwMYG02JIFSfSqRBNL81LPkmX
/knVKpq/pVLHqE8xAI4m/PoyWXnPV+J+I+nnjQPrFkcz0oy4b2S7j8jt1WSeeg6vHgHPTJs105Ac
wl+nH9Lscgq5ytQqOedEvKPfnZEGZqZi4ggeMcdvobcs7ne6e2dRZhMmkCZBnnCYzVvzUbdY8SB0
YXeOMLy8cMd19SvZ5V4Hmj+ZDHS3tngTC/gOnFasDK7gnLa8/0XUIF7W5bJpSCExXxxF2BieZJn7
gWpDceRzfnnAHBjdXexDtPJWZlgAl0T+e349v4eKBLUz64iPbGqtOhddSP+gHn/FayD/NTPk6YlP
JtIPP4aLBWDcH3ofHKqrMZVbZ48qt/zw+s6OPqHKNnFkYSWiV5rkt5s8H1RclCPvsCq+VnhjtUvz
gcaMducScHeqk4W02Ar7Vgz5340CEK55F9zfBFw21OZO9QMROM9qqDneSEbeo6eb663SCJSDF9Ps
fcuQ6vBcSzn17HzOlv3m6GiU7Gvn5m00Fj8XXidgUmjS51kKr62XHb5hEu496Zb6P358KyEq5PVK
UHWfdg8rYURUmtaXRAtdJJvkyLBmbg414yMdQ0Glu/ygJgfeCQfj8y0iL8XSKFM5Cps2ujSjVR20
hltPX+hmB36q13vpUcw3wx354mD11+u84AboDr+7Btp6O0BAOOhX0EMa6Nwb6Y8mHK3/Trjf7zw/
ybVlUG8VdVjowy2NcNOcXcZN4FLL2rK7Jyg+u3GU0c7FKzTmbcqJJak47tsI98BEmvOlEefoRJLt
pIn6epcQ0FWjK3Odwl5vgSxKlqsxicn9DeXa7KkftBRUiy2dCpEuTU1Hh36VF1Xf0OOPPpCagrhC
aZmuchxeadavBFLNBeK1c03MgM0leiZqifLMsCR3Yj2E/f8W/npPGKqW8tx3nRGV4dKyzq/KZ0Cs
Y550+rMQDniFO19NDy7ZvMKEnicDfch6dqbTQoTQWZGVfYMKXF0sRWfmPabzNrUmB2PwFeg7KJA1
rhoPoRJXxJXupvnqsryhvYrOu/99pNdrOzE1eWGUlZtEKmbZcHGSYCWtDbojWUrM2FvVuVOph+/0
3vIl3/fx8OpSBLUieIa8Gd2L2aF4TsLWdILRX7CjYQ1r1K00nv+MZuQndaNxKywufh4wkJMHUTvJ
L6+A55+ZDht2Dxh98tQ3zndae09Rhc6gULr/Mee+NZ/MgJjcBnwvnVu7h5rsPGvRsa/vnD3nXJEr
YGdbNUlIeWORwspxKrcIRSL1mU6ukpkj4Zcaa3DNrE9UOkQKJrh4AFvThVYcmY8M/3JMKHiuFRBz
0gFLHVPAQTN+rf1fuo+O+zqvwSdIqNPCEv+99GlzDfA0ntRC8aMbbsO7doDZRvQ5XERSCjwvSUzr
bF8QYUUFUoERn85Xy6oh10j0mTO44Or+GQFX9c7Tr4smDE5lqqAle+TPyyI3yMWnWaXuJGRmnx3u
hZtQK+6uyx5qoAfpUBq99rBZVOpQABzBN6LxygFoj8+x4G4R7yKlw3Nh+x0ElR41aZd2PkT3o2hU
wJQe5/V4VTLoc/trQ+BhPtD5vT1DLmtklBwr4wC9Z2PfmirMYEAP9Xdeb7rlbtXIdytxr4gf1fyH
txQ0XE2dUtcrCtvJm8p0ioelxxe3Dn0r7xCpUXCiEx3eugFfX5/3KJHnJ7EQQr0fWlUfEtsmksu2
sCwUoiArNLTxIIc1EL+6BOmPV2ltlwWPmDjfKTfBQ68/tymLmpwJxg3tIieKpCMcQ3+HfsO4COsu
NE2BmdWdZM5TWS1PGYomliqMNAzi326jd1eCe8W18TiB9i9WFflc3/1VFgQO74Q3Fs287JEtVBvF
VKsKJEXyFF+L6jPq8TjC7gaBYqY3cwNTb/BxDqdIijmff5xy7oAwlBcP31dZfOVE5cfSlb3BOkUh
yvj0jTji7wCPfz0WJFIKkeNKMkQlVMb/WLup4zRpnqA7E6tk3PI90shlpLt3Ugpk1bjnJkw8cJHN
bFV7kV+tas8o5DbAWTrcO3pdsgUdkqAECBG/X23MS73wN2hwFaFz5tjZNOXHFF7YkhDD/ZDWTiQb
pY7KRlX0NklqsbpN9vy8bP0nHrGO/x1J9nwxfEKZN6vJKxdm+uTgXe+yXPViqYn3KZcuMX30Y3Yv
RJfwAs0M/tx+YGEBfsCQw0XFVauJMXEGX2gF74xN9ybiY7qByh5+FfoWIuXACDkCJvPkBZh8ixv6
9J2dPlq2X/Aq1mzW7FloWK1Pp2jI+R4J10yx/ADYph8786Un4rLJlbY3JyFi8WvqyjJKqZKE6mMT
3sbcuSTLVAtFS1LEu3nECpocQAmZB72hj/g5Q6lTQzSWxMU5wT1ila6mNtVzJBB+ZXOJRGAtfmQw
fo9yL9uw2/SWcvPVbRZ+/9n9inXRd+QlXjj7FP7Qi4W95vtsmH3JrVl8RZ0qoXqB6qWja3ifxWPw
Uz5fThw7wwTs/3ki2rMO32bK2+zByM+yJluzhstpbXUSq/q+FEgXE3QvjOlnmiB88vkpa3M6hLXL
/+o70vhYRDitgUM2zR9sldlEUCk54Ux1eI7JXPDYokeX2S9WeOFgKSfNQn0lqqyy0sqfn3kVO7x4
XKw6L008dXqH3T5uySERLhMW/n1U9YRa2i8eYgOWc/hMz96lZrTGIj4NHwyjULjH5cTmo6M35Ze7
NpHdhOMWvOM/N401PKBBO62LtEKbMnPUKCLW1HIGknItOwpOdE4HOisI3nqz8q7yDWDw9R47Lh6f
iv1C6Iy5rm0oX5w+nOcfxH8LbVAE+2S8n+PVJ+rVowybUxE/jenJWtSDqcaqSFdODBE2tLBz9Zt+
a+eJ+S919Fqv6YSluu0uvEgPt9O60GYY44ITZU2qFhYRZT4e9/3bY+fkUQpdlbObm0oqcJ28avhB
82jxkTfexLnw30eV/9Xspg/8vqkZXoDzhut2ZZueDgwNIPzgJhMmFOVrjpVV5fYEgsCGB6C4gxcZ
4huUw/lUTDV0E6WPv8udh69g+BEowCxVi7KIZwuiKMT+qcjTfTlzWBVACUTHZwixp2iubPVA/G0T
uwBUQtbD6NNzAAvm8k3oiFx3GeA22ccWVfTyrYQ75y1ImzS11BqwQO/hhIUt68X2jb1iK9lQE7Hk
iUyTdtXvurhN5/RQmM3Lay1niXdEJbiHVYa9+AKyGsxYKKTJkmd2WQznC1pZpxRJwHgeHvALdtcF
BeXPelKxypJ6EgpZNJo3IXNOtiLMoW7P1BXznbKB878sRJY5DQ0b5y1aEwleCvmgPXOfRh73Uft7
VFZfdUnR2Wjka9KaWDYGbs0rCKo+h9+jbJMsElp1YfR9OGkeuCNZoS9Cwy7yXECReQejSKQNQzRG
rybrGDH4HTW/JbIi0vmlCMiJOCnnZns8wSCeIePOWdlO1EKP62ZeXxJooHdDEwUzEllF1P5MFlBC
c/tHL57kwQRhaqNSIlDQbu0QkIgv9xV5ud1Hb6uxLNvyfFNiAeI8CLYY2xn9vxKupHgc7RpDlWp9
H2NlG8CBlDGm9C/qeARyi4h1ZN6TsgDL+ocehJIPmYqD4zdgbuiy5EfuIgPm4+rjqOdK+IiT4YDy
sPY6MNjx6r7nvEpqkY59wvAJq18IXxMB8Mn4dPb1ZKW8EKpHL3FwzLq2RGC0TDzD5x1m6W+Nc/6H
CIVfW2gByvZySrOQZVivMMAmyPHHCPYOvBBg6WwSALrGUve6V5+XZWBHI37CLMFs5b9o93Po/yc8
JWvPfhwfF8LHam0P5uu4Oh8R/G3Qj0QXs78jUNwXoynCnTjdn5UD6oDxVpwqiJ0gigl2NAmibmOC
NcDO4sla4LD77C4zmgwSF5vOH4GfhaMbJT+7+F97AfJ+GUOOAT50wD4Uj20wF1H1bVyLQzbqA/zA
F9Y6QC3yBEOua5ivoG8dzzXBkiDqmzIfLVF9mNEmw/sia99sUTJX2zAUSr2o3BJNV6yk871/qCbw
60xElZ+kQtuve10jP31m6LMFoELwc9htaaq2Ue5qJaWRddEICdZJ1utRWMYEf7o60gxn+E9aRcAh
5eBNrLtmJY8Bn68b0ZdaUdEuQCz6ebyqZM/ZiZui4ZnsSLOyBL5CwrrrmiEWL2pszyqXKHZfIUdt
6zd9AgEhq4oLWYlHAo0y4qKfKzFVxs59pVVdp9rCX5MBLJo/ereakGb96xBAWKwmbYmvTNsc74PI
E8K1SRnICIKh3NQQD6g82yH57FwTTeizoylJ5C7f2nzAllyQWFt8xidrTTWg1x3/Uu1OhYYjXNIY
fmnQSFQdoNav1AajM8gcyvnQxaQ7Gpt7bSr4kCyUWh2W8RP2SgOMoM8XI+/yHvOOAYqs2johao6M
iRin0Ka+z7bDpmDKtNBPP7DqOcK13hgG3mn4BMCtmhNud5eyLiYHz/s4uuYWRfeBCFce+H5Dyprt
FcR0v924SOmBxdm6voQAFxPcc7lMIeP76nysWoOe4HbrkQgGRh78qj0C45uN8cU2cXZe9uZRLoDY
G7FkyDy3T4r/SNbwCq+0YApSd+opbWeRj+OUqn2rUyaIAEm7WExMoa9XWVd+YVfL8bteq5jIqtl8
pk/SToTXGYlDH6Os7haQrkdQQuGRrssFhhlhLL+ficc5CIM5oljo67xGXmIrvAVaGM87T0uzYKG+
4Rb26agPCeNpipbfzBQGK2AMJp2hwn8aAL5YTHavdEO6K8W1oEOEr+Lo0aUPsICL+rOJ+1nFLX2s
6dbG4Zn8Y/DN90ZRFncqeXGf/n79T0Vtr/x3bdhyLvsnnHiAX3H74AqY0HJZZCT+ptNL/YoUzMln
izqVCHXOkccc60eV4qQR3sphD/3UM4PiSBGyAMxLBzsfQAQPPtAZGNpWjgInoMH9kLCRdJ+YN0mj
DH2T7h9JeRWgM+pix8Ch6AdPfHYDmBlojObdympISmFRlG7rS4S1Jnf6qmJ37qsY5d1VekSHVxKt
S0Q9WcZQNGxMvNr0o2gXtsP7WpOokPDemXJvo4bTXUszxlfmQncSLJH78kBFSgGUw2OJXW4zlXBA
q2+sH2BFbXoq7Fm1fjFppBmYUKefJuWKmqAAPF3Gsd0QVbARWWlAUxOq/m2zMKaV8iHrnhllz3Ha
1WJZH5eZeB2s/nyO5IiOol+aXbgQPtzDkrBr6S5PDxxs4nqvq0T1nTqQ0YDTgM7dZViCLdPqeYgx
xiADKcO4KQgPdY34vEC75iJTEyjYVLXl5KgSFl5pUKuGTOUID3M/237vnCA7+3KuTi4k3+i4u/Q7
NPNcPLN8Zk6Qky9SV6ecUxuUfrZNBOIYJM+WJo1L+meYZ9oh5DzQ9GOpSS7EZX2S+vTpF8/xJ2Ss
gjZTgBdTAyUIacwS6GXaYn5DfSWPyv2ViseMnV5zq46xe5QvwhJvuaDMVMmmDOSvhoMvxu/kgM4r
Ehesknm7Opcn9x51JI6BQBrt6IvK1wor9gkA1V6l+n3eAGICOtT6NxEb9qs15RwZlMPgWnyv/adD
zn1x3a7OGB1a6/2D6wNuZVrE+eHpTYYg8nx30QvZH/Os7bMDrpwif7v1SMsK/Rl8M7F9ZY2t0/u4
UDoYlQDbDttGjfYTkFySP6EERCo6X+8PhCegR1ue+vZkDATwCQHu+m1BL4J70HvTwYN7SMM1UHYF
Um2vFOHuXq6gN/gCodreCWFKLCQeaYNqe1Dc/8gE0TGjB/utB+2cfFhYLQZsLZh1EIl4ihU4F7Mn
Bd6HBhLdzHNV5ibBHZec/OGZxkcJO8WDCn/aiUo1L70cRwYcGqTRkhMvR2Iw4ia8fxHKdEWpcm7+
LKYdIqP9ff9lsw7EF2zTDTw8Uk3nnyG1Tw0iWlGaTe/N3dqTik/AVwxhNcU6FJ74VrRc3J3SJKQq
1lQgyjfP+sP1d/2QiWQGhx+MLfYPGeiVPhFFhcMkarJVPRmvSS9AGqwiitaJWxa1mk7r9liYFZF0
qzABi7YNtK2zB1jD+KhyCs3nfeCBRKeyPOFVbAEXd3DxO9UlqKtmIZdbe0+m7fSqhGuBiCgdvJKJ
vp1Rzrs7IpZv0FnxFlj2K+0J8/Bb7Rn5upHCfqF2QBmn2OWpT3zF6+q3xB8E1cfnolTjj5xY5zRb
uv4n1sUQIKTK6uobzCnLAAkB9NYeBDN9FxNuSPc85OdCrFJ6moNsaG9S/vm9hRSYI5VNqzLZ/vAa
Z9xpcnyGn8esEetU2izaoeOPVtaOpVyogxqePiSvIR+5/ttSizKpkdOvJ2GT5yKSKIvCd2pHI6YQ
DAXlV8E46K5ek9zzOAxOAbsYHu2WsTtTB7PPnieKm2/dimedQG0ueiT6CmP4B/qBN4zeFsXh2CT2
Iz/2vBtDXhWCgoEb5lfAALz9IMDRIfH2Vo6KsPZtYvi9wfKWR65x5fZmOEYAsmOPMJp9E/Eb2ELw
ufLzPKT+/AUu1C8kKGlWBimhRW968mXbn1Yzpljwtks6LDx1Wb48BJC7BDC5YS31alZtOCek+cm+
VOL6J47nol/DzPRRHKbMLswzmQchWf5PPgeZstfKG5w4cGfUON98SNruAlHiN3jmaefaFdOo4q5F
GLZmWXJZxFr1Lb3KpjVDqZTZF20I+Osnw+yqgLsX+8GvSu9rqYoQGBclSdFUak99uaxr75d8ie3Z
58Lbr1GXvMd4vB7teZBlxY3aw8Bjtc8sCdHlV/eyWT8e6rHqZ1zS+RMB4EOFbA4zeTX5b/AqU6w8
+J5bPZCS14EJ/Ynj63eM+4jTHDawvyE7phNd3ZUJ3nBuCbw37XjsWonUSderIMZlXTia1Tb+R9a/
yDpWQRu24E9WiGQGiwclNU/alXLOY6F0xW/4Ybp+YN4HGPYFxP5vAhBEwn+pQsYMyHNUw7gXqXOR
C0roAsDLdJolHNcDeCea7GvpEYwtdxLvg0W+LS5R7lgwd5uwJIoUPDrwrX7gHVpDJ9lXFmwsYabw
3I/qU1ODVV0ZQztJbxaIPQP9LujQlnuvOWsftUqkM87nJNokczkJGvTkC+LpOE/rjEcLE3C7OQs4
HIl4GNic3Sim1VlmTK0At4V0gx7rPMuJPNNInSayXZy/AxhqAUNaO/YQbxc1s1bvw0YAqrEadStP
f1p+iGPo0fUtaB2azxmMVbL47ZwdSp40jig4Z5+WHCiVEIV1de6w4rGaUpfQSwb96JEyLCUW/ZQ/
5UbIxBIbDPwUXLY3pmUTOaG0aVZ2AGwMLsG0fzhW4kwVJnBrdswRb4u+qr9fmj9wQjUDmFFoLRgf
NCo4O4PPAPdS1DuVycebkPppMf9d4zceXGeM3fXKML1Vss9MHwPUjhTXGFVuG0tKxBflKQD+ETnE
tA+CbTk8mqAa2drgvz3Yn9WVaUUq0d5kFqgwowf02j/zpMeMFzyraf85ffiHvF+qU8uq5/ie2X+m
C3pGHhgsZZQZ6Vwdxj0oAoalKzLqIm9r1fReGuDhk6GtOlndH4x0iuPCD4VlCl1dNM/ccOPpJ6Ad
d2MK774gPHW8K737GTzvJDQQQIUBnlvpNQEVWAwS4nLSHdjW3CfHgWPJ4YEchBCS6yS5zMtS3A5S
GpalxQCB2x88F5DlgjPqfO5RLBlK2ySyGWTScpoQgsSoNaIC8Qs6su/SN+I5k6GnqbDbaTtA11wl
dEKmeSJiZ4XbSKKxgiKdH0/3Aq8c4vPKQ+GdWtKpck09lVWw6l40jAjw87ajWhli4q6psDFroGif
u2aC8myIX7/FzWLw6lQzzpDs8t26tngxbCEKCxgddFpVPFsAryACo4iE8IUAa6mnr/vFNPYajTl7
0O3fjI8+JkqYUW3irdX+OZPVFopSmNAZWuMEDjHLwC3ng0dRey8x1ZfXgYNvZjIc1wwD140fa+bc
yGy+6N0wP+DQsKSpUv3HSGzGoCD5Ex5C8d59iXcmeW9TXRJH2/KadjlUOO4iTzX1Nfrvf5ccXM1f
cbpZ574MT+69TQP24mNCWTJRR85ADQw06pDcNpq+2fJvXRxk21dWkc4zeI2VFPY/XWiq3NNUm0kt
MzOFzLd9+D53CdHpP0a9Bv6u/GABdU8VPsFjtjZ2vRhzXCs8UTDNSx6yeSRk7/8F0Jik1sj+06Ix
otLA2tz8bRpFElA5yyAhiHIaa7pXzbzhQaYOAq9gSAnZQrGZPfphNwI8oZXw8V+hrDbuWPW6BfiT
UAJ0hnLtxnKxWjZNrIimMGDXqYG52eudP2mbZ51HPuZIXMU94mYUUTxKcxNj4RqoJn2EYCjeEwht
HwNbRbmsxnSwh3zasXqSXYL9ugcrQBBe3XQfgafr7rPGpydAzC0iRlgy1TRN81CaaYLB8tTIH5aq
wFTYInC0MFGqKgKAKF1LKdFwz6Jp7H0m5unAWSxvIhzcfbs0db1MiZBlrp/u2CWVrZyMSsX5jaub
yiz9sPl+5qKvu3RtmsCVfk7pQOGzHqwh7cgpCEpO5/G8blBMhE0QsT0/uUdkK+yQBme8mN6OPOp7
8K3vJaYoBx/Rd4UjW36X9oukmbweNM4TqnH7aHutk2TbdMb2P5Bb0aQT4TYHv9TnPQ2I5MA4xcZf
CBUp3Gjuu9SxmPggVuUuUBmp0H9CQ+i3Di0ynS5x/Yw1ufoJFksLe7u/t3GsWt+CXf9LtE4qPd8u
sBiCpXF1JbMu/lCrDZ8j7TZDiXVt6PEHSTUJLsJK3U6sUBecx2PGTfdklgL79nqKdEuBkw1HWYSt
qJvcSGosaCN9MyzYh+CgLh4BWAPsTaNChdXlIlEWVWbhEopI5WCJiOBc56nO2WyNQmy/lF0xDRVX
l7H4zanPMlyJfqspSBQfKzQPbrvGOY87ReL6N3g2hEkaxYNGKujTUVmgsHEOE+Q35ZgDfcvMKHD8
r1L9+RcTxHxTB0KbtIGgofbJDVGbvOFmD0bRZn4JwZXOupUZ8CerdtwHKfXLEnQAgwuuwAYb1C2m
OrTviFGkr/4+TvG30lndixnXrjLqdC6eu+jmuahaTE8PEYu1PiBcD+fy72Y84W9+4SAu9k8HRFnu
Pgc9azacgARJGmbRtyPDo9gqEd9FDhhRKqwtNM55bRcLyLPFij7uFUWjcCF7bIiSajJgvOsN0SGA
zsAY9++pSJxzhdMZP4UbbzwhzLRy4IjwJrMf/ygY5JqeCHGnISvTSK3eTDBVgKBKImoyf+6xy5ji
5KuSX22fHv9xpjOaY+9iQsISuKaFi+2hBkOiVfzUXCq15Knoa54CIToCmHYqmuERyGdZObVFKzm6
cNPSfCHWQ4wXnOYRfAU2q9pezdBAckQOzjRTRvluLG3M6E+1II8BDVma8SrNzXJwfHXmxea0T82q
E7lQNswXMqqpCh2Acy/Asg96wDOewuEcOD5nRHthH2xPJ5z9tqO0gCsG3QM7uALBJTa3DCbZyUVg
KX/QdLTrdCRasJ527Jx/X0/Ky9amdKMJPQypG8Fa837Yyf9McbPnJGCNCCMZ/EEfmE/taRbtpXo0
fkX/Qlfxx3TniAk7Rb/hKXhMOWTthCLBYbaZVdUt4da47QM6Saapyzzq9Y/0dBz8BIHGoIPEAFwr
R0MhS7PFtANn1QBCe8WwAu5zobr2nSF5/nbiUjefVWpx6qaFBNlV2QeRlcKpzsNNcAsRxoqLk7e2
CChulwDhUlk2u6CrqCU6ZIyR6lhS/CaypAr4r3jZCU8L4RrsokFMq6Fh0wL8cpEvUovl7c5V4teJ
OkV56cPNXle1/nQ7+o/5eAmfPV/igczvxOXDOpkGy3WQ0bqJP1lm1jbLboZWIrALIFerU9f+yPc9
T5ObHIFww65kz/6m5KJElbnzDw1EcmNQ0IxUr23cti15855jhxeGKqB9O60U3aRxt6kKMa5IEnxa
C3xhKGbGdaqsS9l4XjLHaUgOQzWj0QiUr+QO4G/K3/UGHQR0ZNH7beP4s/1b5RelZQDCaraZBRak
I4p7mCOQ8dP+sYnSvlPLTlKrWCAW6yHF6bhd5YMwOSM1TQOGRPycZL7gs/HrWyomk0/rv2XAi2vt
Aw5lDdv6ufYuX6ycuVY2zVRocmIcIbzPzRcNyMydyNCVHrKPs5qgfqWPPnkmHp8FBUyrMVPr1pfc
RAeWQKBmUB9beJSX/0Fb80sZCCwbGK+aAv36DeI1Z2SVnacwO/yYbjN6j/wLZockhIyouPktGZUt
YfQ6OwbcA5G5e6c0M1QK/0LEPXnEjxxENsDsQtRBfpHVpEEF8g2Pf2D0Qa5aOX2Y2jbVcTRG6oVi
hda8lYV6pJmiDGKiAnca1eIhqbxaftaOG5uW73eSXjuywoRCfx4NHbuRqGnddxY5RyTA7zj4Ccu7
15fb9IVtz0T09OWgVtcKuwMBXW9hXUFxfUSUASxkXWTACVPLEsyMz5ExfIfV2hOoNirfpibH9aSk
Rh7yTWQpmlQwvdZNchHqOBuWAhrulcT8aKWP15QIe86Do9APsxm57cm2uUooxhFS2tsSeR+dcuWn
xBtN+ANLpAjZMrdS+pNqi+6MOtTKvRewdJUziWv6ER3B6Rhl4IzdiA8hh+lYTN7UlPVEkIDmxz+H
Aq5AQRivRjaenJvIRYhQzUzBNgFpujNFIMgUooEz4lt5U3cFT6HeIKQW/fRIox8noA5gj+4YphD9
QuhSX7qhhTeSaoYhvPDwAOyRFRImp+k+cmwdWkyvjxlVbkHT8ZuVGnOarqeZeVZJDfWGiGowYZl8
3X2icv/COEOqMSkNvs56qWr2+U1qnVZoeqIKUNBQQfvIShUgcMkHOaYvHBikgej6LLqFrF2HHX54
RBt/ElnlsL0atiTF7zWzkEXbAWRfxfwE6uf33YSmpCm2c3coLU2AJvHjE4Jb+knM7NMPj+JavDqX
9vyipMcj/f88KD530RYmPhYd5M1NIEo5B5SGHa8Pf4VYlvQJOtNfNjNsORZhnO+2aXAObe0JK9mW
ob7WArFfOiYGvbyaDgLM+qmnBGDv2hiL2nrsLIjp91NBg0+kL4qTfzsphzrwc/ii5U57kn8dISv9
LeQl7pBkV8ugBtHK+dnj8k6Be0I8hbS13WVZ0PtWmcROiZOBsUAcbQB5SVVnH4V0oeXWum4Qcefg
fb9dEMlebZd65nyQSSa1YOpDbplJmDdEFvIvIRzDE+hVoGcQSWY0+IO/8eZAnGDKqUXNlcDIN72p
zVFERGCV/OiF1wFZOt/evptGAFGPGjB8voM1hVQPzLn0UpgxhFi2rWmY+YAwTLUYBt/X1pTyQwvF
KiM3dX/6IU/QxP+/u1SpCX3QQyHvMqkfKY3Qt6Y9clkgemIkg7X0ERCqKIu5T5CEojw3skNZFeVM
IeIME985PQUe/v0XX7yJVGxRKALHzSKW0A2Uw7gM9zXXbsAOAsIlm/daq9xytZm2T3kP8wgulXfy
MY6Qd27Zmse+RzQqSzMkeDXeG7dVAwA3+i/Nr3R+TGp+WE7ZeHcbCUVTq6WjNU8PtkvFwAvmynrE
St8KTsLuXTC3283r4r7eX5P4WO/971j252h2Bz9o2gBlS/NBphzqnJCsJMA+csAvpEfYaDEE4Nr2
kOOKa1xHKUcxR1RpLojrBWuj4uX6D0I5N7Wn5kKgz0Y1Jc9tn0LUnJZzzX64IxgKW9UV5J++ZBlI
vW9qDYX3pCmjfgEIRgIemzilCSM2Ao+aGVeAX+q1WWEbVHjz3trUYwPwUyyEM5MPLhwW0UzXHI8J
w+b+JgXcm6BiMSwO1OnqmDq5naPq43hQ5wSROaX09eUVQpyG8xs2pBok4xTnB2B7QlRsY3PYKFO5
G0l9cM5qeVK37p+KcireggW+kp4u7+sTmEEsYCAcc+8+aax3RvB6zhSNmpDfUYUK5kwYQHUHwRiB
qjuI8PfoBNBuv45cBL4kpwJO1wvRkQg3lqeu/c8Kwt3NskPA8YF5ngTbW9TJudIEquDoyBRmpC86
2ivryhaBnKT+xpEYOF9eZYoXjVelkUx0Md0spluZ0cyXDfAo0HQv5NdYA47HjncowgUhPqKZEQXv
TNFe6tLb1xxg++b+J8T1N0d3LkNDAsasMWqSibMTOVfz7PERirB2SEDN3vWn9SuDSsxBrPmEktQt
oZE+mfEnyHTs0IAyE3s8bxABeTM5CGylUSkFudVOZp7ZqiEUGP7e9vAfGsDzWs1giouFuhBbJ5go
UVY9aC49wGw700yx4UciNzFiWDUN0LHgoZJX3QTWm/bowtEiWmeF6KbokiqYnIg+u0LfeMFOFUwy
Ek4LrjRoKPsRqt3YnrhHR4jQXd8HWqILV1z+fyibEyCr9HVi7/r+NAHyLLPWVeYjq+231rApkrNS
x6I+Qp9mNwDNjYP4FaJbqqUDaZEUSB8tZNtICJ4pxe728s/XNy3XYLMvxQHJe5d6VfE/tCiaUBvU
g5f2pAg1i1I4yKyx8GefwImoaFP3/KO9kZ2lWPGhue+ZStUj3ig/+qSNSrIJwm9mgZ5O6pDRDHi3
O6Xg8auPrN316m9I8V9D6f9jvxTG1LClGpu+byVZ5NO5k5J58h5jF0KzhFUOrbRooqmnQ+1IpUyh
R9wB7PFx/BFLiRTljaR3KrETdishYmNkeVSqKPFgMCw03Gf3+fIcQMhg89C8hF7O29BhkMYWf1SI
1DBPb7DtEYVgCQHetknFbid47rBxNxRvtm8WpRM2jqAjEkgjy/qFFoBP6onqlu7aqTwDBhu6iL58
cQ40qF34eqEKoRglrGO9M5YjRzH/Izu2XmPQrk74rwaDTvMsDWGCCAg9gfMTqbKhsLI1uRAD7hLA
1rSXkFtazLE5qCg01bWMDlcp7nZlpd0olZI7sAGJOQrIbFGaIQ4LQ3pM2f6NBpjfnzR5/ss1tUwC
8wNrHekHarpBnTDvr1RFEXjvyjKVOsSdGu3vVOWX3hS2btXXjCgjVF7HNxxPki2S0TW/zII2v/Mj
3aXo5Rdk/ZhkJv3xWvRIK4V15VEtF5455iiZYAfGdKmQVqdU9+nOHts9ynrOvcmV0npv0U1qO+F1
Zn7ihelFriCSe+yomXnUZt9+xq0f3p20vURBQdEhO4BW15FrpVurt53Hg0U47lWUGmJroF7J05rD
4+x0oSs0tr+CkyWkYK3x4c6bpZqb/d2XE7p+sZw8m7vtFlcyTl5eO1bUVb13UNAJc/l07uRpJTbN
D1nRrBRuD5gWaa2XSW+S4A/PdZ6ZHkWeMh7SH4G8KLvKxpA8SpoY+8hQwGcLR1b4LeRK3MWyHOxg
M+9sFaM6mAh0hg/7qQoxETCLKpcvRycOcq32vtcf3jBHulht+q1dCzVKo6lfzZxQ3SjgcYIEOVMX
l/mSMq+p5bXXM3fYorXyIV923O8ozb/XsePiLu/KJqg5dDqfmCS3nKecJJEcBQBsyIf0Z+CYBjNe
se7noY5v1shH/w+GuhQbHARSxmIKJM1d6I8r6A05CeamfymB4HiAPYRJKq0ZFlnfRaOOiN/2m4Dq
N6q45gH9xvpChflp/ayPrNuUmBeXdvsgLeLFH2dBVVQg3AlZGcRxgYUrRZxrvPCXosbT3zpBZTcf
qznlMeyKbB18LoyMh6tocU+O5QyfTQHvT3W46WTFK887EfvYLv8HEYTveBCwUZ54Eu/EpbJiq3Y2
PfnBc7WTSgGH+4tcifoClsaMazpJMyBX3ePr9J1dW+8OtXCBIzEgcGT0fweBDr8RPO/fGWZdr5C+
PY6eB1teNW4ihkKbXEk1G3ZBwzSwbe+msvgaSLTpWLKCRI3hUmnzqKLnQmsXYLRg7H+eLiP7to3K
UZLL5xz1pcOMc3ABcKeovr5J0W9v4rgvu+gr6gA3d3XBp25dr/5yObM6h5S5S/9HxYJQBEGcJPGv
VWjW+RD+JLG5CT2OxyIK6TOJz6w/6ocbGm3E8sRSYGs18FWGEMix+EvzfnUGr2Bi9lnKLP7RWOt1
50ymg0XVJUSBHtyYvp7DjBZYuP5uFI8D1EENuY1YTbWjsQihBd8P/acp0ciM0zf58c5U/aCH3aQ1
JSQfyGjag/+DUNEnQlx9dIt6UCu932SZDeB29g1iFmIOxHDEv483WBkFjp/ocnQKoG5HSP1Xuhoc
IoWgaGwSLXuw/j66z5zbM176xm+YYGSXi5nkgvFm8Zqj1D82wwhquJ/bPzrRmSHd+aKW4UbqtJXb
TT+JwbpZvhW9fClDKFfZspOESnjskCC0FalPPinrHo68WPXwmjfnAxAVHzh0aGgviWu6GJ/vrz+Y
V0tKChEWi5sZm3hF6VQ1zU9f/ple0j8W7r090o3NX/2sz5l4G63UulWn+Ui6YDq0gA2qI+5otUwG
j4kOWe6YQU0H+kKTHH8bydpaUcaOIMlH3l5+sKCLCcQr/GvDhTwjunGUEJa0xIIVLembGCD/YySC
XUjDtZfeIG9FLD5dg3XFjIIVwmZa82anyvo5qOS5izwMCU4Tb1HbKg8iE7WnCwZZUdYnVdgxSdbR
X+ZG3nNa1NEHf+wJ3mEf2DEJYwLSUArh7NsaGlfnSG9Vaw4fbVotvLgp5l+jUk8QKN6iZCf/SGu9
vPupDa9WnD3yAwEkE1DzQriY2Mc2N/qjm0eo+6jtdRghejMgH1ySxKnwciaTyokSPlr5Xj0VEJTU
xMC3KGn0GuoArtp0PHjPL/f5q90qfYwZ5pw7DeLoW1kSniV3xhG0HkZV0E7n36/pUx+tO7qJXs5f
nA3MDHgSFdTIka/rYK5Cifvz/t7vssRaPxVnU0L3EWtXXsSzGXWx2rMGrM2rDVqOoFJyGH1uXw2P
+zcpjQ2Iytn7c2VBPvRukU9oL4cDS/dmHNEh9hblPdfrGeyAnrwOulFDG899kGRp/9oFrOkCmWMB
mjJhhAdhy5VNCNvZaaqkTCjNUweIVuUdqAXGwZoUtMr1R2IkXTQNxjx8+ji0Nzp7pknbAm1hv80Q
H8vAHFv8lWqSPHDMPifR2R/YBumOt9OiwYtMmLfi2v9quQlXgfcwdRA4LkSflw9Ob887OCjscvf5
Aan4LSwcZrvqYYTNSu8XZJ2dWYNkNpeuefNvZKljMAUhutj4TBPy/Sr3IPWM21FTXAJ17ivTZSK0
tvthE/1ZfgyMh7N2gvFZTKOo0AJB1HBaZZUFChFZNU203sBWU8aTOUPImo+SPtAixLBtesmqBcx+
nOuaIQzvwmjuD4QcG1kbElrMbQKxn05nN0vzW1b/wMDhp0XiL9d5MEKyXQpR6wUSx632PMqGy/uZ
MbvLi15csm4bhGwDWFBk8xBS6iGXtm302TeUk5EmdxQW21NiphoGxJkW7By1FVAtjoOuiYtwJ8sQ
pKJS/HQBbz4kQbAHwr6an68QooSj26zaAq0hzEsIS/9/ySvPnunW1NkB4xeobkiteGPh5ltLu9cz
gUGIQavAvzKEJzyyrraRuJDneAJw4wGY2fK7FOFN5PiIzfKBZaWEnDSwfUz/hrWi2r6H2imdY2FZ
cpbN+DCcQm/IoVRVhk3/fQVAJVcOogpuJMuvbNVmCtVt5cilc0FRCsvqWFC+07AGi4XOu6u4Ar2n
l8LN7cTCs7L+jVc0OtVQXbOaRMRqaY19QWj4rCzwdUmg0Ad0sJQ9H/db3COYINYT8c7LaKT0k8EE
58mwxslLn+aVghUWKOwD+zl4ww+NgAXWLt2tysI4l9+tsDAGmDYH1tFlYj/sqXFVNl5H7Yl1Chzb
T5BTS8nS6yH7CrQD23hEzlJesYMT6Dc1ewqRhooWXmDeowONQEhXGOMdvJmOsRXaaprLsqouMjoJ
ZvzgXoSZYyXmecQckgIDzcaE7G7iYM1Ldh3ysWB2RGiDrKuXJ8IiaLWxsOIHNSI6iAKo6UQxVgYF
1NdrOq3WvaPWeYMfiRa2aU4ovnKtFNpTuS1AS95BCQF8BwiEBrZca4UV/JQIJbcG+pEZ3KfD/gxo
4jB7RYA4Q9IL9GCb5XBp6s0Bjb7slnDqU9Gruxv2i+Y7BMUCVnF2KC7aXOjs2U1jBmN1K4UoIbog
BsibBhvNun0K+aL4gtxsR+xWTMiCyaDQsLbrTsuDu+81xB4EU2GOUq7C2hG7G8j+Ov3QonUbG+Ab
psjXRPzHK07/JvsZX10DWPFFzLEkfzcQua9x3uO/bX9timQFmCn++AY/vGIQu3htta+1D1yWqEBU
aJno1WUnkys5K3rAtMn1qWcn+O/GO3UhEmedpAX4pgPxlTSe0RJT3Lm5UZXRiyc9QFlx8noUDTSQ
TDaEDCUILpPgVwVubCbv+p38B5bw5hicqt4ADoNwXV7YvCL//Bn25h3itUXM3zYjn/84nzBFhA0m
8uWRNmhe0rAUOFiMieG+RnnpuL08A7RczPABUdsLx0iA5QIKiB1hgyXs4oSBHvvGyFDyAH7yVfRF
C07L+G/Z4n57lJ73+AyR0SxwWfTdmYxFut4OorFc2kD4UHvGOsDD/EnIS1usUxjHS+/9wTt+waF9
oUbApSEw2s0AU+h+6eH/D8wc2oxlxD2LC07LkUlh9nArc1p+79yhRldbGB5cF7B9YEEhiNU4mQlK
zPZ/iWql3KZu2BWM+ou+f+IPZKDC3csVp0N5340T4QX8UQ4wTLYgTTa/Dm5Xp/nKdvxCTo7D5Pgs
oQpBjdhZEwfJD1xPp0+hbAtx5swQwqmuT7doLsv+CFUFI6A/+Sspl206RyIEIF8WcfyNVj5RnUGJ
/oKD7/lBF679AIXGi7OZAR4LqufLe62Vb3X/cJOl7Yc6mdcxXfhyIdJVdHyRsLN5S6zbyz3iLUcr
oD8oogIza1wpGfNxPOQF4yBlrlENFnyZt5ApVKVPE3D6RBP/Pk77F6QahvryDoY9ZRzckb0t+b7Z
Vv80TYbnYNmlktENopXMkwH1M360Y7vDbg+HQMpDqC21vTg4EXM9g+bzr5Rh1tCkYI9Puk/gTo9E
/zyPZFsITT87YaMeYkVGZ1XlszNH7fbb5PNmqwAlX47cGC8nDSw1m7XSDbP3V97IKy9U80s3v/Ad
UJ1NtG1CxGj3fpgvjLu+zmd/Xua4S7UWrLFoub5i65oMhfsmPMhlhksLrd9AMeWPgvMTWCOCEiok
7O/EaRR3rrXqJQ9Njl8RzhA1fMGx9zB+p0tErZh3FEsW4ZN38NyDH0SjtvYvo4fEWpAdftKPhg8H
l1EQH+XxB3pyOVYkYotv5dKRnLTAWQHucUztCM15AOetdJSBBqn13RY/pg6VC8/D3F5sbv9Vlms6
9jTMSDDOuks2EbyX/snBli4sjmlOeKUhX16b5lRoz7yIJ3mCm8rCTsBxOwz/OB//p8V9/Q3moKcn
Av9+Fp1IIhpcSzawSiNcS36gfu/2n8+R+Ug6ZByA3NF582ywMgHly8HfJ+Cwj711jDCJMfwx7mo2
55VoRAiyBu27V31jlOK8NxpXeVIiu7paKt9M586fuvrCWsVEuFufoOxAKTZdwO9prq0KFWRGiOI8
NFlAzMSPSVIREqaIwXzLD831vnfQ15hllXu5hzLKX4YhoTtYrE/XXg7b7ctDE6XiGwQq6mXoJE3h
VxVj7gMrLCBGqGdfm4i9gitV6MJHlLLt261ewuUobXR3OvEfXoe/CGf4HdjQGx6siCur/ERV4+4P
SuPRLhHbd+hLqLbYdq8yWyjvLoKakcV8Ez/8OdqQdeFhcobX8X8wksWvwM73DehKCmpf3VVIYK4d
YH/PGwd0qruJwTvCfydH0Ss7EbFFA2VsUiSkwvBySBZlWD+1cE4AxPrzUozWc1TPK8Eb6zRu2GiL
437ug1i8/TmFhPGVfUGu+OAKkhg2U8kDlONE8u2HvlG/Gkgjf8ZQA3ICW0uiY0WXMC0pfkGaM+33
asqpZCaMzYo74O8dA5yaaPBRJKD+5uaag08vMLiH18Yyisw/1Bl46AdsyZJCA8rt1qCUFPXwYos8
d6A5loB7iqxspDKFq7lnLWa6DxBUT3xC1EHOmIVCuuLBJOjZ5NUeoExX15yzmClIKL5qBlkAgOpg
rFeUoo++0ZA6FdeqhFigJcPL3LaxSWyCzp3aI41As1RuX4Nrv8V+dcskIInlk+jV0aV/nRdrFujE
RaaDgeMHmKOVRvK9r1ggGmJvfX+q2x081JfjfgoRVhNeZU8dIb5Ibj0DnHj4KYJsrBPy+PbQnwn9
6mj9RZBf7KClnc5wXBGLM2460mNmmIT/i4EvVEgIQ2BLQ/9RxCnTyxwhuj5GN22aXWl+5MrbZanX
iDCRySK9H/75k5kKOHCd3s+CpetLTKN3Tpeq5/kRlgGjk6NvSKpe5FptcrnsvoD1XCTkINRvnYbd
hOnNIafnmeymxippWZxVf02aQ/i/Btw8ffg0B7BywmZ42Ej4f7lhozOddq+GE5L13vjVmM3cEkOE
QfcM+6dtm7NaWk5oAGq89uDKK4VMz4TkuxInle782rz38AgN2RE4y4uvSD0TgCXesn4lUJqA6c07
IDPFPpy8fprNf1HFxpTHWixGEKOJwSljiJ6MH5aEK3WTkfdm5kSICo8FW2d4eJSOCBFtb+DaQGw8
u8jfTMwdANv8BxPKnpepow/4AGufznFPCEfupNc7wysPuYck8PcMxWpIxLRorqjbq5c3KvSvh1sI
hHEYZBgXrLKHYJIUQO/J5IjOI9LFielHUqT6w7BhIrVFp7pvCn6+ksJEH+jeRinxhEf6V40EXOlg
utzzyQMDS4tONtXvI80UhxgaDewfNOsx8p+jpQfshUH05NjqA5JFaHYS+HcI9ku29avLQhdVP6MN
VniSQh4uNFfhY7K1vosAZrw551lHcGX+iuvOqaGeKl9bNFQ2kxWi3Pq5DAZvoymrqrXZolPXsAWh
jprfnHz3ji7iLvXo4wYULbVdWtjHvkPCQ99KRtkfzlqBiztk1VfIf6rQBFFppj+6ijZWStfvtYDK
7KsaflZ0Z9EBLmuws4m+ZoDBA2zXzq35UExohH88wMYh6Nt85G7LWmeMBJDwvWh/QiTSkRmBPiiV
99cwJMMdMYazJCNfUjB2Lq4FDZEWcVp1EiA351b5kiifVppU26tZ74f6LJHgejyUoTIuq9bNwjIf
As8owt12N44/cJKiiekiZEznCR1wG9GF93A89lIe2wf2RcvLql+Q2OwCHrpkAkQDOgTD7gFdCqpa
0uSGc3/bdOPiysC1QJ+XTNLkH7/UCFxMAz8PgpLlqfdTZVbZY7DB16gSrAGZVhHVrBpWZnUAXBLW
8qGUC1yBxsvyj3uvo76kDP0acF2OyJWLYRhUsanq9pcdSI60JhaWj3Sap3SqOVFyyGoCr/OY2Ol8
D6fBM9lFZ03gztf+8LjNp0qVLFE8G6vzuVgcuC5IHEOs4F9MOm5RXMi6AOqoQlZ5zcZKxgQ0L8h8
kYhZMxxKvlbZ8KXuzRtU76G8/lToZ3acM3rRQcJU5bPWkcRRN1GfXVk+AljQostCZDcbndfUjWDB
2KFiXOcsjZD2LQ+YUPTSsuyfYhwhozVM/ryvpl3/rZAqI/7k9WMHGQPYQoOgNwLFqxRew+ohmzKd
rmX54w14U5lTw/IZYRcYTfg9xmMzT9oXKKxEie8XcHmYbtjvnJ5+WYuMbz/5q0S591leAkNxGkPs
2mir4o1dzSTsWTeuoHXmSQ1/RGeXNoL7sbse84/w1cW7abTpKVORZTGhhR8vRll5FF1QTBQ7iNV+
vVeymSJvTkENCzwd2O02R3lhqTJi7xmsFgGtzNkt9sKOL3K9/TrNnLyBiZzwbtg87fcNyINEVH4R
XaNzCH4cn9fV3lRB/fGEXPKuJgrahZjrGrfiksiF2bc3r2Iy7P7QVDpSkWmeMcZKp8fAfnShj4JK
DlBa+TejMM61BRRUVJEGzHlWx3CoNsINHELyWKlAw/eyYlfnzjCTn0GBfLxzUAcs/QDkZXfrSDUB
5znLxExytds4TryFm+hWN0yg+fFTHLEk22tMoCEIBCuSgSmgvb6/xRKRGxSyoDYE8Gpe0BZQWi9e
9ph6SxrGCw1Ew5zCJ/l5bRazhlS4xw7MGrVApuPqpfumYEIUJDILBOpvMGQZK9WiGpeSSlPimiyV
8Ww2RpifqAt/Ixa0CazhybVUqboBQj7N1Xgax1guDE7nJAnECqxAFrZ81kySUArKcbH/TO1ZKDBo
E65RZEJXqZhilvJyTL8H00i3WH6mFp27pEKROOEDfYVsdJEDG+C0TK0v15VxnuKTLlazGySToZpw
sgItSSYVGUT0Q39lcVlaY9IWLom6zAANYyn5mS5VPplsO5tuEwF0xrYNlTj5AmD11clRrXHu1n5+
lYTrpk3ROK9B7qXYeVjrjLHCTL85GsZ966dH5pVRqZadVIN4gHZZkXlS0iAyhm/MhVX1HHk18gh/
wz/vOIeRmwGAe5ev/RF3izNymuo7qcrQdCJhNkmGagwhnk3hjYBsd7N+ZAzl92sw0UdFpfPU6N5Z
yo8wlFkkAXgUmn46gFUL7gJlGk8QUR9J3LPV53jG2/NkquvxVX5G+jiTTg/lxgrvb54AaKO+H8BR
o/uPdDM+wund9CM79Bc/S2Cn5Bqv21pZU1M/WR6kW4wQWe+XRWzdupWDgjZrCHCOBz0cIH1j71Ru
Xj8j8j4if8QrTZYJragt79Ws9wKPhufbbx0zOn0FWB3Ob7oyk/TIBc7w2rgNzdnC1gklB4ML2BYr
yvjBbK8XjV9sso4DgahW2ICS6r90U4PzAEobjyesjXXQ1tYYOqhVWv4bHEdh9L5YYc6rQdmFtOCt
myPwgkLk6T3ob7kBGFet5FKW/cxAzCi11CNsG3InvySHKyCv6Hh2bfV2jhslLU/UOvtWt5XKLLo2
3fAE3QYXCcVlNLXxYeHX5BjqWrYUrAB6xmmlQbxZyBOI9va5ZhmBCY//XxCOzTTATHWNsFjnhzXx
FK0+OCGMoWtmDamhwQ15UZbtRATCGM4ZIDFzoJtPqsNnHNEeC+lkyoB+rjUtcBUjCIr12oGK2MIO
aIoD0lbj/TIqx6kD/CKgj1UlRxT4Wv41cS/cSsKKE/iW3ung1KrEfUiP/076RIDXnSDvREnWgp0f
1+st6Hao/mzgMtB/FKKJzkJCuek39iXrhmzh6AoTCzUBPc2T/GVMotY6DN8o+A9wwIkEXha8K8n7
D4Y+4rg88zFlAP1GaZIICBkZ+CFLKkqCaagTYOgiOWrCMZoq3FshUIVvnQ5/w28D7HkA5Lfy3EmQ
QtrghAi034a25YcEClou997fBwcPhaRQRHHD3GP3T5oOtiGRUHmXOnugx43xLEdCLjT6/2C9vXN1
piYuNTjF3bIDawOr0nSFzS5XDCJyveAvW3XpkfIYMdLIoH9uI8q0y1+LHlLYmMapf8UspU5dUWUh
XPiLuu6gqgG9Nl1sZ9EDctwdmyqfEGw3yrf48Kr9OzACdnmi0JgbP2LPWr6EID/z1+uwIFglz1QG
d9mSX692UQ02dgHtyF/mBrmzAfvwSdJMARJjGsDmfHJUtp996tKHZosOmIIeb6Oww7fzoS9zx3CB
WJbW9iZ3quSE4957mqGZpohdawRBiGt25TNAEWVu4RjvDMOiqf8jfFjDnUb/kA8CEAIzHjoSGFj4
172D8g/xD61SXg5+ClFlC1AQAV2hlDVY3dI3ReNtMY3E7fccqU5atEBCpHfikC0Uq+9Xp6xLV1Zq
gyGiCERLraKbWMX4wB+LN/cYTpfJ6FF+QLqVY6WGYjk4QgsZmkk9JVWSYbB5yCYDdeiAh+1JkLLP
8lom0Ue20bKCXgnPUlSroQld224+SJV87qZv4L6mXMvMOjY5izpqoKj7kZ47nBdGMZCLK9Dm0RO/
WeiWwIQbeZbxlEbPM5rPkAJ36jjSJHvSRcsT0C4YnWy9vWGSmB8njs9sbfL0Ihe5H6+rFsUc3Uj7
UQ5i9PRYHVEAhKOJAGHMHGFHcgBB0MnDAfoRIrsf1INs414yI6uQQKJH0Nmk0+gpLW1RYMOlBdfJ
LGmdKisQvYebkxJ7ycRqVNdc2QDp3pDbripJc809dYlGEfFdDomuJ0rFp/337odwOBVTQNp5ucd5
MgL5BVKaAF9wxirTXwPmFWFthaDUN+Kz6cZJbv5+5ZVoYD6zSnKYyh+wLkWVaRseOD6pc3ylHHNr
4QMoFiJrK/rW3bg9t9RlFS2zuNvoRubn7RFHIwFBwrDQjLhZpA0AwrPgZM1sjhxKR6XGPwG4L2/2
945XjQcHMsKTxEAbGhILhuJrDxYgSNLz8hjJoxxYQ8z14hrtdVofyGCZfrpjZEvN5Xje8p3qImGM
CVlAqyJ3zm84WizkwjAgH6iELXYiYvwqPnDiT9RctnBHeFDUgUjgj/zJ9pqHwrAwZ/cgHRtLWOgX
TDECFOPtGRo/3l9syzXIZ3LPH0qnO8OR1RUIoTh5uD709ARgl8NjPHl//z3IXlIcyPxZpdrt5Lag
HFQdzni6Dw4uHkgRjb3tB3sOhnhHcqFJkafKHGyNuwgZbZWqa/17ZWCJSKivIcIW9B8XecUyXtLh
bh0P0U5l16DUvVFSVIHjFRB03fxkSLqTV+xxpInTy8TgLqER7PyGy359IAMeoeJJyZCmBJ6FjguW
aOWldh28hlSd4bvG+GZtJyBe3FW6T8N54YmnOmw07smPOWER1JmOXZtmiDTC1e1CxUDIqjYCpdIx
D52WIjis2Bek1V6EpX2i2YgqvWnSTZ1g2UgvnAzfh5uDJ/Mp5UwGxcFs8YF7IJ4Jha6P78rl8hda
I/LbDdMdNW7rr4eWh996R3Tfg8MkEPOL0/DI8/Zn0sEFOETDglv0KbDpU1e8iIaSwOyFU+j0RP5p
pyFppv/IeZ7acAOydhWT/kAxWJl16Ri4NJ9dqSaHX/icBG1vhPWKfM0kXVBbyv5hHyRu/Vh6pvb/
vQpgpXK75ACUTehh35PHQFxJmSbZSLOHvuMD98w7SLrORehYkyRUpqF9fLrwPxKQwc0gf7VtvQxu
PnzXNmYU4xFR7mSN9AUWIkUZDiAvp6mAAkdoaNUsxsXQd8/Xf8NwXQbmDew9o/epMHqDfNXb3CiV
s3xQYNurfwdMJhcx3LaAf3np2BD2nNPInLrn6GxeLCdybpzwr92eIomzyhg5ONpx0eMJzg4DqHoK
cZdephKovsSVSbEJ/u9MvjiGceder6xqZk5aDE8v5l824KCm3hiHXroan0gx4IPl5tKbG7l7n9wa
Mcpf+GUii+TJsAL3CSjouQXz7AEj3lZJ3AzUGj56wravlpXUfuskR6iP0teh8TdEMBqyfVOh7iqS
t7ZlPIvXyYDCnNJwB+QaRY0xikeNBgT1vLqI677fenBWUrCeggkZVMWZ1ustZcfjvX8Yi63pMgmS
HFY8RHv1RDc5DIjwQpLeQo7nWdaCA3j+8aq8AjZJBAkKeHUwY++j1GEQLzPdlBNzi0NO3z57X/3l
zrLMcNZMOroD4jK2vDfzf9+M4BAAoGI6uAI/kfHI8tzuX4E7z9FI5EcwFBEgGFnhHxtRqMgCmM1+
5S+F+CI6zA5rJO1FISZ0YknIVyip7JWHcCjBNu1e5+TcI6wXVzNmb9gA6dqQtcnKj5K1NK1J8HvS
7StTK6vzt88fmB9JqMBeKsfxH2PTnvspPJabdhHdYuH9tF58RveNu4HMK6O+qUd+2nEg6+LwG7dH
JqJGzpwYtJcYjhU2xDQBXmD36M/NbabZjJfvwD3ck+6D3W3PY6LHMGLDgSvT6l6KykYtTiMo1ia+
W0LABezOxf1yxooPGZrEMRSD34hUSb2GvrETob/bU6AuR7YK3FcfP8x4vpSegeMcGfPJ8pgXJtfb
lI/UxeY8c07u7dLyuahJPNgA+fiAHRb5NBB33oL/H2e/eSl8INrD/KZrQmKzey2cWZ35kKuB1Ws1
AxYuc6F/6r+741epW4iQcwjnhXgPq3W09Y1HVTP0L3ZqGRLFIGh4Mu7YmtUfATuM2zjM79CUP03f
uIRgQh5SnGJq4Kb9MvMMZ1Fx6kK4cDP3ayJWGJDq06PCavZ+XvuG5T+D+6hfec79w6xkUllAn3kL
iPZQlMpWpNAh8Oq5QwylyyA1PRAf/OqnFTbKO+2vQmokeNQ7qdCwLs1Ssy3WMvQIxD2zYHBjxWb0
woiwvWmmzwEZKu6IFvINVsOAn2EF2VUMfezc0dw+pgLNX1lYGU42hts6AnAV1n8XaoEVMj5lelm+
zh83msNRVesmSMVZXAYTTHnuNQkLjFQOaIIZzBVHUQLbvzojYoUxfWCdS/Kb7G9xmrI/G2YF/eZw
/DIl7yqfM3UWBjM6Gi0bcUR0bjQYMBwWczuwVoVVkWj6jW1/EimgRCHC/sTwigyC96BrGZxOwN8f
/M3G0xBW9jJKr0noRCzmMqaCLiocgcY05eNBXAt0IZRLBAVQix1ijwCT6KGntORENYjR+uGARafw
F1gnrf6QUPIDZ8YHnp3pEuPMeKDt/K65Q5fsrCOOkJ0vjIvISPSxFhMAZcPS9o5mp8e9CD41B54S
vP7tvpqiiCRrjB+BXZa+nAlVF+ubrsMiczf0c/Jf/BVRrx7stcamwhPta6IMbJQxryVXb49k8OJI
5mN2DruYen2FJ5mbtSA57VaGKBI5PkOA/yxrwdmfbx7Ls6FLBNbJCpsMEt2u+rMbuw/ty4AXBIPb
1PlwwNnGfmPQPlS8EDponc53u+E4KBsOIk2pmyak34GI305IPZGt3zrWeHy1WQxdN2TdgH52V1ao
UTXecSLdd478sloS9Za4IzJH9unormwuqCnXY7RAc7qzavhrYvJysOCyqm8QWeO2D/miyk8jBD1T
Zj5sZMqe5YjeVFUkIiFlmHa8ym+3/8QjusBmRRu8HySMd65b4UBW+LVyHFoPW+dEMnjT00JFCoUo
iA1u8jb211RCs+rCqm+wvNaWLnjSFdtnoaBDt+Rtcyy4KNV27/JGBO3ZyyI0AVgy/kzKTjrGHFaL
l2td0NQqRaNbn7H3Kt2QeO7btwUxfYf/cuyYdaAprY1ltfuWElh34ubkfsdU48V7AWLFxJQnOO8F
iYtRCmZGCkdjfLbcaoBS3mMWaeKPmsWCZPS2B9ZJehUTugCb1T7Ui0gsS5i/cExI6ILJM2tNdmZz
8zh0jv7fM8iGmiahQ3pdArmbHnh1Iv0xR9BbsbPMl1yn8gzTbCix4aGJEIUz5PcU3h1HeFpkA5TX
U0iUDJqLejgPiFPxHcvcdSvnHj5Bt9hq1bMJmM+2LhEGp90gCBpOtSnEQsGakTXxycl74/iCdQcF
QJO0L4jLVszedpTqQE3MgGzpGUDb84mSL2cXqVFo8Kibf9o0VzPuSG4MpWMPhQvCy3augYDKYEe1
52K5xVeFUPqZJgIyG2aGLWTC5hK0s7wCCYEgOHsIBlxrnB19xjW6WSkdEdOghW0Ict+BEoOr4Eq1
hV+u4pZoMYe3Jj7T6f4GmfOitR3aa03MFQXUF2EzpeGZGZwk8EhSBGTuBJwxvuOFfgAjX7WIc8ev
zW4L4n2Ao3jdTsDuM6yBnzF8z6cDUaqbPfwwlEH5L/3iMopF7GINXXP2NsgNTk7d9oSkR3GXMWcF
RDchPMu68cBTB5ZT3GOC2QT2r7cEFA3yrMV4OVzbmOlemhqNG/lMWrgP6Pvu77q5n6JS51pma9Y0
4eCxlsKQt8m1XGOFiDrQm2jfuOdiRchB8lOyM34T6fMbGctbQq9Q5ukO3deP+mO4LaAVh2SEIcxO
OCCa6VUJcZ04X7Psm/ZHQ+KjuFpFu1dUkxRQKHuw42NLrpTwfc7YAGLcuiYIJtztXZ6zJZq3TACQ
KK7RX5PrMHCXOz2oP2r+wSsBFj2Xys4LoNLdJ+gCq5mmLYoIV0aJ2S9hRQWAovS3T7iKnRlPth51
jIhdQHvHWTtZZpNf+8SWpvTvzBbSn2+ymkP2zouHZlQJbG16PJch4m2JxlKpCZXRIYEqLAC96vaJ
9fHgG/nj4j5Fe5X9/7KRy0+AI3bY03thbOS8CG9Z0TjzqhXNdjXlmZbRMAZfM8P6pFKt5jqs26UM
10g6oYk9P8GMZQj2BNfjFQgV4TTw6xT6mRLy35obyR6eDFbQEYl9EF3w8G4/sJ9aneSwooDyr9R8
Qcf2+LDsjAJfpykaXyW1R3ldShjZz+FsPdnbyebTU1/QCB35UJz7HfFKXHbgku6R04rxKRyz1GH2
DWKiurP3Bz8tjF7EWCzlSA0an9zD0vFruAQEiFr6i6/0IwIn8z4PUJR4O2oIImZbAW8CJFBFGiyp
NXHR/RreUfp3+o8cYzrm9Wum5e3Ps2MmSRUdgJ6Y/r5LYk9xDjLlRzGtSrpx1cOZN3n1lYn9qAw2
gzGZhnYZlTDJU5AH4RPGSgqvL16SgxBgbdgUji/BfdnAkZSGoRX4wjjrWeaAP525O0os7B91ONPm
pOZSQTIkI9GJZJqkSn/rNCofRuOyADeJhf8A4mxtZ85e9xrYinhwqZXiR1UUba0F6iV6ObkhdFAT
5TcrQzbyqEK35h9W1R/C1HgXrmzCuGlRbDH16P7zo+XQhakDwl46zgqEKxPbF/1sWa8h5qqevU3I
/7ORWguyP63U6M8mirajpQ9G6wY1XuDDtzKZZo2DThSOhqU3GWJPUB/ITFxcmqDIiRYtOV+qn3Xg
Y719FXxAeqCeMO1qdbGH72mlr3uj9Znu8Ru/W7SB6WREyFdYL701Cod9xeM2cgT9keNHQ3bI7tff
Ln+QfYFnLxh1v5X8lerjPDu4AqvKM6S9LORw0Zn2xeEFzAFM9WoZo/QtPOfUNQiZKzyOW/PHX680
BP2p1ozegmSbNTuJJjp+BL4UugmhX2wWQjSslYOpZe41kplF+wGE7qvk+3lgy1DY7QUne+BB5gpi
nA1p3DyD3d5qUZ3GmvgZ57HLtSOLc8Qkfcwm/No1H9mtxNpmfiDPleZhiVsEUvio3TXCiU1uit5M
mzVBPRYW3uqInoXyOjHHgMe0de+BD7XLmkDwNrXTOmPFBmLL64yc8dP8uveaghlrL/2oSJmN3Nek
k39cWTMn3KHezhI1Pg4oZ9UHj47VR72/gWAYXdofGlYHqhpESjw7oCRrdzO1+krzDM4YMfWU+WYZ
5+CEDerP28MfHcPq1ILf3aOXedRAL/B9FzPHVVw1uKkBtj8B0kmpBxC967LQQBQCxBU6Eu19qnkR
nvHUyUCafGrv2/HCVzTu+itEu+av0lk1Tdq+ZNL3ZuBgnutzGthaCkYLn4bmcp3q/q6mi4LCNJZl
JDfJaRDOvtWIsOrR9FAybx9zanqT7a3tvXFa2OhjA6ZQnD5fQB3BQPw//7eyqepkgoo/rfieD3Jj
CXANWDTtlUJWbO8hM985WRJPGkvtZg32wMRLT2E1lhq5K2g+pZFJ1wFY3j7bDQ4KrM+rPXYGYfsM
IeEoRME+VZaa7zX0f7Z21fMXkUVXNo3y8V+FOnLb1OshZ8auqCMNObDsOo2mIBNe3QKBTfi86YTF
isfLPH7QSQfz0tyRx8bUWm58heMomOjVkfIQYVoRlocdwB8+gouQt+A9Tkn+zUICzxUPqkUKkUln
SKyLsQp3VJ6Es9N1Sigo5ly6PDqAXGz9O/8Fy0Farz4uW8u3vuj+qjSbKpETyNuVY29OnA827+BA
sHGZ72M4c7VPXGvguIKQQJF89SzdAsxKNJOn5qezlnpAHezVZW1zW6a9XT/Ub9GACr8VAIMh1c5f
VV2VzPghQPH7+zJuQrCrGUE4Ojp4aNAToNV0hBhGfzYIcUfCofnaxp0Yyb/oXu5spwX0B6E3wXAB
3ft15Tv21IFAc9XlxLuzP6jB92Ntsvynafl/cbzzNR4tZTxTYXgumhFE5EMWDyeugogaMfQbDpo1
Acy1KaxEyew3JVFllcj3WfCFOrCNyGYtZZDrcULCDYoRDeAvw5DTYlS6F5EH8zl3gzj7Z1D9r4kp
8X7MzsZPQCQ8+i/IjDNoo+pYSOaok34l1OgOfGGfz6hJAUCcreMXTqr3fhBIpD8bj7Lzt791W2ui
wrLjLlsDueZnmaGl4q31PSfoEM2/28pCMjP1Th4jlb9WOy60bT42YC1fRe3YDTXKLAuFQxlWC4JZ
QTg/DVjHSlJzuxSOTW8dpYIe+2lejrI/jJdkHNrc2fIZIB2mdXDV5RhT6lpbCYrIC3S5+ijXfZav
7t6mvPNJg4FkVyCplBt63PXEag2soI+Kbuieqxt4ZibMvmZlQZYRF+qaqJNLYoZwJlUad8afK/RR
2vv3+NNWKeSiPDBYQxnYXTyJo5mExTEQIgRtTNZTiBsSKepPiOqQvt7dne4A2WRyVSaZ2PcI86XM
E0fQkPQZfif70vmGu3qZMwmMBxoZgoirTz3OA2MOVqQDTksh82NuhYsJJw79Cjm8CLJjPEizyH0h
9aSq8IHHb+ygKssPZ06SCJ7prGa5awTurcuWScZSzUniPVk0JdAjQfP7yPtP8mj+xaiQqx61udHU
FPY0eAdi8AgDbne+8kbfb2Nwxik6OuAZQAuCxskupqmfB0QgHqlfdsRgnNf18V2pMNEly4Zz4q5F
Ke29RYoER5lCe6CGXSmxp1/iZzjMb2gxU7KcoL0YFpfnUZ6cbxhHGnr8bLmHHACj3AnmTiDWWYXs
joru8fEkjBHpBADusCUiaB8s2jmQtYA9Z3FPNGFMRGjDydAgDeT95wSfwzZ25LjS/wCUHBe6SEzv
0GDZKKMoobVbWtabnkt9Nh4qzmyvda/V/SNUmQMXr9iRXMoNh7lHly2C/jtlCr+P4KIfpLcyAzh2
90BPgLGXMCg9KrhFXMzUBj3gIASJJKsFhOHxd08qFxnsyRJcLlDy/qqmzGgX8cm/BSC5bUBAhCq7
oItCuN1bIZoMry5V2KMTuNtqIVrh9cNdXQA5GBYYB2gDKFEMkEA5qrscEyT1Jm0tmx0u+2sgjR37
upyG8rQHWNYwLlshKUt3q6iOfmi8A/UyxJLPzQOXdFt33D+yB5fYUY53jqDZmmpaq2LjuKEj0zs3
OdYy5rAdOzY1bjYg0tHqDBuf17YGl6i6p+3Q9WraLQPklJgcM/p+0/lUvduTvwvb+Y1Ybthdow4A
oWj4ofggS0/OBQ4jLwa+WFxqDlFbnC+8V89JO3EI45WFabSsXrVN+wF+IuCFH2f4dMUE6jl7YcBQ
9Ka4j+5h0lK6l1sE9XScyAT4VNFi2D3BQU8wIsaRlRmPOSfsmfJUjHDlhumfLMuRzbysauDkCP/C
WwawPF7h4JLCc5BeMqC4Itvv5s4gGbhac1/Q7tkH0TUbPY2mhwQhMRk0BHwmpnf0A3qP2FqPeo5G
Y7sHe0xoBDMT8Gqqa3DebudY8kEn439ljlIqjmFtwGx1XgGsIqePHusgqkVtSIvo3nPFN9AZcYjl
aMOXU1GuRtUrY20ubHVz6fUgI8HhjQMkpFuqjq4/XrzsuGOnSqnfkKm6meQiZgOQMTkdRfFrau5+
KjJbmTOCKXvc8FOnxfq+FPAx48Lzq6PmkmQ5x1I0dzExTr2xUHlmDYjH2d+A9LgwRKi2ZxoMiGzf
XkB0S6tn9rKMzoSKO5zo8mt9QkkOrKT6ilRjkf6rOFPNtk/WAvShwEB2Gc6jQQeTFNoH5LOc7yiD
B6RtYBlQCj3IbnSFNQdSolIRKo3O5Mb8jKLPUqesaO875w+lFdd29ljD/MUKAyf5RpqMgKbkAm73
rqDf9k1CuKi/fNRk+cqbrOGR+5/XQY2luDqbnMYxAvRDY0LNyNH1AEJ+HmHj+zyseNku+pfaztzF
c9CXtwPWnJw1pTh+DrHUkUxkRxVOjN0UlRjCAU8X/8vG6cgbRp4i2zXnU/Exjbc84ZWFSZTMn0I5
w9Wgu/x8WavOIgJUnRc4MdWqmVB146LhBi+erkk4z8Kz6GL5T3/cbiwyIk0RSHIl38CH5u91MBvk
gftCu5n5Rz31Lsjts8JOJJhJTiFGYUNy7rmLr0LnQXEj4fMUZSd5fRmtR0zVgsyUg7Aql3AmLfUW
e/zAXp1XFk4LfIaxc1ifvGWqjaE2/YZ4J7zgMmYYjZd11o5AzTOnuXkCfPLTcIbjA5R6F5id625w
ZJ6FvJD7VceDvyMjFzJxWFhqvF5qlZ9b3gVYUa71NHIuCfZQF7qzm2f3P2L+WWq/IKTeTIx6IWje
Y51Z1XO8YmGjkrE9Hja7FyTwXX3O9EQhej6tYZXGECWYiZ/m33lMkael2aN30gXD+CAXtiighC7H
nsIlkZM/FLq1iXKj0snex5Ic/cJDdl2H9gBCSkoPJOz9niIFJhfY3Upg9Qv/kt0IrXAyZxWtXtRX
wlZlLA13/KHu0TkMtWlOGdiC+u/znKFMyxIIoBliLMFOyFyo0FWVE6ZBEW04y32RgnugeJGhLvf1
hzTDeZlchu9iyRIiPSeEbt/chWHHT5pFef1a90wpV73QGWxRxgiBpzkQzzbKzndsBG5gfSpEFH8c
HVaoUa7Ev3Xv70p6cp8eESbNbSScEapQgE1qyHy69DHu2UjXyB3Un9QQcoDfmsZ0uLKV93sEKCcF
aCG52C/o5BHh8ZvnWpt84LDSDzAFXu6O50GMRtIoR629NgQvhvmXhWcIlCEdMh+b89qcTFwF0tTE
DN5T8FWbcOw0D5iKXlZPAIlUR4Cm3Y8/8QAIvB0BiPNtWCMIeJ2r7gpT1J84GpFaGDktanz7Hszn
uVVekvyeOVCIIrtTZ2GokwbSS+oP7E31atRuEUfs3GC6JLldmHKuC++No0fguY3FREMeVljanez7
a6AJr17ZmRgjw7Eoks9hYQGzuqAVX6EzIH+JrfkKFXGQxcB0YVvOiOkryDSXkLMYclgEPdgTwHVx
iKtJgpwrJFC2JXiOe8wCNKiGS9yzcDA8Hnkufg8DlB6HoyddESdEXpLm1TapsLbKoADDwRVGQEVo
BB0Ls8OULX9UukZ974VRJi2fQYh47uh08ksjW4cvUYI8Ih67zPqXtC+q6meeakIfpVv7wps246sD
S5qyG9GREXTgRQkL2bjZTIvkLctcaVjwwT5ol1qNR4HDOqTCYqlixw1/JjVYkFelqajtQqWaHS8C
jFd3R4LJalXW8iBotCaODzVE1UmVPoAIDg5jrD4d8bWZi4/EN4o5ScbHDNZHD+8WjPBb/QBRQ+tu
XaYtNE4t9m8o2tRwRdHLS3xam9o8evSQSTGnCXMTsKvd4y7gGH6LGAJ3aDYE1p/4LodysmtoTZNv
NsmUDjeORYuyUOul+U1fFIP0Xom6q8hxSZuO3a4QhEc4zt1cbe9hJEwPpjdnGV/oZuI1920ofvhz
pkJ0NTxhkUUwlgQGWQTP81eNXvf2IqeHi1uq9/+8pJ48eu5jGkXxTzM6Y0LEwauichJ8dqSXVBdx
sbWzf81MNdIg21j5TTqjWwm4jmwH+kk5zxtkVNKGLB40VWoaqfbJhy8Io7lvfn+6wf2NxkvT8YQt
XUz6b5EoKLkZVXJmryUDd/i1ilfAlhQ7gCHpnaqhWNlX1xmBnimci+bDWlVzP4Bz0CwSPDnIbBXl
j54WxXtBXkjZmKMGGjNlLu8GAZ6gJo8hOsAPmkxIuK9bcw9hPfatJqB1z4pAAuqjqXbdEY5Qyzqx
SSKcRiIh4LXxDnEFFBuT4yBbTB7WNzLr9H+73CNqvOwNatBF2FRLV90AeNLXI8Jnd3I3ClgWbHWa
JbjXn4Q139vkTyrfJU/EyDlOElx0WxCFQ52wudDO1F0qT8SDdav/Bh4E4YhuiYV7QE1TUvWXNNpG
GHNlasHesjLocnzuVhe34Zw9GIPVz8cC6Fg2i3mzUaVZu5BQE7vHmr4ujtYHhj8u/BL85XEVdYsc
5x3Rn/2XXOJOW5lT+bIKLJehr1NdxXlh1WuHOZ+xvxXS7DpALrL6ldL6QflYCKcBEG9uEycpkAAC
sIl7JwVu6BTf8hTKfsI4ZaHJSUg6Eryrtdcg0TNYAhLTk0/BnCCQDx6Xlb3dr+IovBohxTy6DNcQ
fLELFBgOAsX2fcwhqQDgV3b1J8y4gbihk6sk9wGc61tgUW2qihtI2b143eyeYPrRuuk+6zJ7eIzt
M8dmagOY2rlpkmv+YwspiF92x8ExkG75bx6/+aHnnQMuciiH/uDUnusU90K9zltD1o4uVYOuMhDD
60WS23UvnQL/kpzB0Gw6j12x0DnIxBSMdjI9yIQ+j9oqIGHHK32Inab7ZMKS5G6OTpFVA/CGjb0M
qEIUtlQEPXDOsrPywnDn0pyfWPVyZiAtbr1IkA1kFsJSaxVs3Vld4X4UYPENQgnyOuUYDW3XaPVk
IUGNFg1LFszf5GGnN8zoYHU5n/S9rHoCpPTU7jfH/U2A2EKTJxLswfadRxJKYB/jtk0BwXUShqkZ
/w69p5PtTof9TcYzJKAR4NJvVjbXC7VOTlDL8zQBKoMb/6Ih/J1yaBF2bOEpTtLhKBrkmYBm5K/x
1rKL2qWynsVMdjgo2PogRWRR+zvIPQsBvAs8yk5tiSzMDp9TIdVlQYX0qb0zvlRLu0z3dYkTtC94
oEPsbtvzxxU2OFwlGagpD/amSHgv9wXdNctrsRZqSPk8ZYasQgjMw310aJv6Nwg5HR0oaZKQOOSQ
zjJQOyZOonkYdFXHy5cQrO+Ipvxcst8OaOl6RzVBYZ/xoi583FJQML0DVywAY0V73mJJhDdUKtnT
ZTK9k7/5efGFH1Uz3+w26SkbDJul0H98c60uP9bLyx4ZNbqvNnDyCXGSCIeq9VFUgqihGhvnWsQO
iqSPF9Z1b4aU38JkS1WndOQHavveDOvfOHb0mOZFGc+iCjfTWF8SCvZ7XuRqgDnoUimyQUENYEto
UJYWPGG4EPicfNm+5c3VljXz71q7IhuxIfu4oCMlaNkiSbXpcIL88otGwBYk341P2mJbYCDSRJMC
xNjqLUZKuHyyCvQLW/6E4siBVp9GoknUm6j28Rpn34qD1vXO9rP4STajO0TXeW7Tk9biinIM7sUJ
mC0KyEAZ/AsBTm3VYpd9crxzA/dXQzT14BE/phcrKPRloij10cE8w8zihSLmOfx4k+L3MrxTpaB0
IKIO/sSoK+WYOanBL85okL6PLQiuON/O4asnv2tmiahps0DClPIEhdhYGMwqWRDDrPrGd61XLaS+
TGjPyi7z9w7YFiKGxSPWbs9M0AXgCeaIS0H/mpMBDp8NLC8H0JazWaqZgkNDuYQiaqXy+MCCxo8r
u/cPLC22okv0E6+ALBeRxZNtcyZRHdQLkwxK50+cUSx499UWGTHkOfcPlVNUHcCIH4VQQ7d1cqSe
fDecXOWalhboxMk9ewUiIEhaE82NDHz2sDMFxw3hg6Ig1P5M2ePw0tGZGyfCWk1YFf+w//7Q9w8Q
Rrs1VdK0faWEKLWUQX5AiiCooKdYUCNvyqnOfoVCUn8sT1XmxD+CsMHMxpT76/p8sQdq5Yot76rY
xwLM2AshIhmq4H/ZaQMLyNp8sSkmMntVXkfFXEqVYlM5wMp4BGLVNTwiiPWEMJlwrWyFeYpM50SB
HSohH1iB3L3OJrE2crbOIfcqICz02u4PDRRXfbBpFweTcVbiHJ7ym8FhqRzhFYjWCnerruGvo66D
6CG98gkI09hPbiNcNgxB/Sg5hhL0ZAsMepLBmuAo0SDtsLgFOdwSdBNNReAIs5SK/S6kIUQ7Cl3W
EJHaTg2A/Zc1VY+w0zXcu8vflSxUxSTM1mrEwzVrUP5QZiGSKRS6kf0jonqR060IosHHRYGX3Cr6
+VN97sgC4z/aG/wLdwDDoO6p3Lx9kMtMKKMaKJDJWAvgPv/Pm2c67f74aInm2Y+39l44KGl4QaD6
mWo3U0OSIZ++eM5yKhebLPA56zBRHxTnPzkBhyCl6xNCXycUIjYab+tvg1VCYuf4d0u7ihu6knmN
CUFUkolonsLdf2nkMm82w9aSsiKyYa0bMpDkT8R9Tkw+PdHRYS4vq707jzHAx/s9pqzj7kL0x7SS
2/2fG8TWMfIYBufT0SPP9ZpJpaC1EkzPq89FMpmzMDkNHi6RhZ6ecsnFOzW7Sq7ukUAHLI8NwZZh
g1QDg6RaB7xukmXGqrf5+u5y2jcSyWgfJMliFwsUF9TznKtUnqt1CRy4deQ/Q9MRRduLrl5wJ4/p
gyrtpQahV3B4/9dfb515rI7uXwfXGuw5pskCFInxMgTm02jLAYecPU1RgjmtiWKYbyPUivpkSBEU
AV/mx5ATHCMwcZnjeFSMYPEpb3+Gyzwa3iiXDCXmn697fkH+S9AxYfbblB1nwCRQXYPqcHMgMlw5
Fa0D2Utcr5gVaJS9Q+HgqRuW9nxAyUaup991mx1Nb90C+cYARtwQqeZ0wFNOoFfKwCqDfiqvzQnE
ps9b41tnRbrgQXgEzRRIaqF3SWuZr6i7svQZDMesS+pii+yYT9yiKHJBvOifCt6aC3nhRsSkmcT6
aHkiN9Dwdr+QSNMcyO479x/UV2DM3O6ZbJeH/v8TOolrvNA4TyM1wzEmCVI3me8ELLf2znX+UpMa
YTkDRBkS0WgMBHk3KEnabcOA0sN8O7SFpQTYMYQYv3TUX9G390Z8OUx7XR+Yy/yLWpbC2Jmaf1ft
0slbLHnM/b5+tMD0WD3wQ02jCRevhM7U7Ai6m66a6QmvV847DCP1PnUivUvY84vYQ7Cv/jxslkoW
2Cg5mki+45G57xUUwTDbGlf1ZkGNEyHDO79Uf/raJwtTmi/WLGUehvIcCFn93SJOEXTzqZK6LGPl
ODTgdyUb1tvfobtUDVj2z2EIVaxb+V8ALHoCywHEr2OFXgLwWv4Wx6qqYCdlVKMfUdt4x5iJtytz
Y2uDFnhELx4kpdPXxLJ0mt8eEqiYEnKoXAk+Al5xzrwgYxnQkXPqRm0JsEs793c3jPoHLII3tKT+
Y31KN0aihFqrXppeOv5gNVq0svNoiJx51aqtnHnj5E0AzJWEis8WKi+M7/DawKjLf3gC6c7WyL3r
Jd4lUxTd44ctSlNltTT7D1qshSB8x4Fqgl3vXcAjQgz8JBaqR+oC2Sk3KifCGtlmDwehKu8scB1a
QMn8DJjdprp4SRUdkiEoGYLAoajOkkcgaduMlCQBt1pApgU/DyY2K75BNS/AynaVKjOkdHswj9Ii
9m73VHBjlmtHFI2ST72ItzzNLVhvERlBCunJOQrtGcjqHt4IBzZ2OpmQjucKKKHQydLn5Jo91YPW
aZECoymYbcmgRSkm+1OUth4MjcKoXr9R7ZpPzwtHLWlfylfN/AWJjTToJKJXpRcACf44brDwTq40
d5VRwBUwtFJdSd13tqmTPuti3q4g0NhFHrVsOLdPRPcNaqCTj1BV5gluWzQWvQS6WU1zfYpZ3U9g
jOt+ab61i+4t5oZZuev//95SxwJq5mab6oYy4JJ9QZkYO0xjUhlWg+RKxSzf1XRN8qKw0nd/oZ1n
sXrUgruOkMiEmWDxOOsxqm3XHCDLbSSWQvRs6HuegIz53gAs0Dreatrx6Mt4DRpvZno4apQ83TfB
p1jpVfhwZNy9A/QFSRCn/IHD4rTnrpTEN0N7h03OPLTp9ANTgqOvL+VYLqrbIKRse7SNO7HfzhWa
ZLeDrcL2lramYG5bAZBRx81Of2ZLDVrzEfHSNOMNL6lOxQS2ncNRmZGRG/y2fC5reNoWI1RZYL4V
eVXPfr5jpcirnAAL2gu2Mebaofn+84yyx3p/NrFtBa488gS02NcSPNBTUtvFpicEqdo1j9Iz4KI2
jj91xgmva9KbEK4VdDlzwygoNExL5OpQ8EF9EIFL/4rATAYI5FccL5QmyVFTliueELLNC8ysKiP3
oSrcY/aKc3W6iVkCAAs7VczO3vqWYGWqHcCZmgcEM7kycCeWimFR5n6G6igavm3rwGbY9GmsOodN
W79zXHWPosQ/EeI41gW9fUflDOYFfGzCuErXrwr6w5vRCWHcTYDu0/c2oiHqlfevb8HwQR816XZ+
jF3pOzatiKGeOxCctUpdjsJG6eB5pnCfkRtvtsYtS/vIbNl0KuQmKvVnt5S3HWHVnYAq4dMZRdcI
8KVQeq5qYkYZtHX5UG7o0UEczlYYOCxRunQhhbiwpLMJz9YcrpX4KKxHF1bc0405j6jL0aykaoGV
ac7hMlgpk/cS/s0pJ0vjdpKmbsuyNaXPRzG1HHUccWwT1hxMPG2lf1Os9X6csMlDEuynznYmYoec
YUAEKPG6Co2XEeLAlVd+I8znaj+plbeO1LaPRomB25CRJRzcWRfc4SpoW/pQkhzINK7JmYTzt9t6
Cjpei3qLCCSFSOtaDl5z4AKE6q0he7AqZi8B+teDhluXKwTV2yob5B6z9AUE4X1Ep+ixq6uVaBxk
Zzl+Aqs2bruMm8zD+ZbwUCWrGEomTg15SyM+iaHnMbzrszCnFFfQNM/IT1kbsGmmlkXIYMwYGGse
fb/5HHCIeKSEsEWdg0vV0sIqme1JJt7nL9AeoZVIxDoDuYFrJtzC2AvwK+XS9lraE/grPIyl5qoR
15nw55JBXGK7XasQT2zcpMhWR+ZjnsXZ9fbnZHv6pa72iEUWH/YmaJhMqe9Cks9tKdbgqCnuJyfn
JUVtwW22S86cgXqdO+Srd5sUGJ29WCGEMiNypbLGPUJO2gI146jCz80uBORo4MmC/YxV2SvkQ5b0
+RoomRZnHPbtGQrVHfoRIVfZvTxXPsykTzLZRxRfXFqN4GGlWDNn67DYk+0dW8CMmjkzFbfbEwOk
YvL9n3lx/IfupgtCunitq+CI0DzyGbIhTj1LumrPGov13GRNO2jVM8gYcQTUDXa4Tu6Vt9oUr8nQ
AS73v4WfU+MbS2WJiiTSunu6c6Mcg/QdiUmI0BzmMD7SsA0sBp0G2DdnS1f9FVCD7x5QiNCL+hiz
iBhJgCKkHV0GxZteI4rAxUAAW1iWAAGMpT8wc0yWjqPuTqanEo+0mvrte6hKNKW+CUspiHkcRVu5
0wzNQulkXmiIJ47OxJZGqQAwC2Hb8XSe+6tXdNcu4qDDEZrZQAl/KOHOjKc3Qzv5cfZSH/xAWn/0
ZUnzdCJBoS7S1RDUaaNPYPWcYc6IpHsYt/mG5rLR3jY3Og0dzKEM8Ba2duW3WW/Cero++EUWUF2t
k8nE92fpDWsugnJVr9sDXiM11lwlQp33mLj3g2u8ZUDCp1Y3bBy5hmT9sWP4giZ8iAX88K4oM5L0
11FeZZtlrcf3vItx1VkCWTIs7u56MVaHg4JQmnZDkU+atOrAZEpkvOzQ0hY+eLK7iQzETaftTbQd
U+NTMbDctuvPwoI16aNFT2Yk+kLhmoraYxjh6HAAj9CyQo22cXprbQB0NTElCN7Z/tCHRKM/Wj+d
oCm3vQGe4rbjYjbJRhUjfn2oJz1MIzVzzt2MdSgq74zIcTuomrBv/yvaUrNidzH9+6puv+iXH6yN
lMNF95VTBkS0M+yYj/FRWON1xW1IXvYj17C9l+ffaa5yvoCLvHqloHcWopJp44WLTC0xUor+6TdC
OckCtlyVVhBGF/A619QEDYQ9gtfdJDypXCl9Q+ooTKCy3m3BaQH/Ottg6ABzu3yjDE7lOONwVRc0
bd4Ok5I5rIkknPAdMav1bI9wVavUip2Sg8RpYkUzl1LGl8fsI+/TR5k4hHAorW2obkA4vpWQRInQ
flMMGT/G0LnX1445QVnxHX2IhGVX04WbqH12hKznCMW5tAvqtkrX7fvcXmYQ/tXhStcwaljoU/Vi
bwekqLxipDaaxoy2QkcC+s7jq+IMj2v21FRhXQhoewU5VuqboW1mRtvA+yjQcf6CiDb5B6fMnyNR
CsZbIhQ2MoJwgiQNiya1/G7zuTLF3SdFMDP0u8JqWiBXOErHuGEU0RRL7n0Uny6mCs/uMM6fyeM3
BwsWCV8FedDkAh3dR5UHxS+0pnODvCBzA6cRaoGSEVj2gD+Zh2AMkgCdz7bXrOSrc7HJRuIQLr8/
Ht7pdyR90nRiCUV5YF77e9UJAvNHwhHyCsyFxZzMjg25+nf9fkU6WkiK9Qj6oEybqzkfHXyRI/ou
0tBr7m0V2MHViyw3BKlohwRclB0hEHcTpNJZlgNzIO6JZhlfGMZDNzStaVy+YRk/V5I+X93dfcU6
E/YeM6N++im1xTgvLyGXOU0cx5dasZrki13BBWAMRn9RfiGhgyVyM/8zEI6QCyfq4AIGlr0IodrS
jIypp93PYNSLc9rtw1DllBpd12S8rGtBMPJqK+8jqQSIxK2iama5z/liNFWxDTtl7xW8hxppvfMb
rbU/LwSfM9bS+pEp2xyIG12wc5Ue1qTmc63wDs036K++g3GFRmo6ChH17R4SeiI9LWB8wCCJSzXQ
u3IkMGcWHjPScZU0sdaRIdSSuhYbCZ4hQXyr7s1xDu03va/9LDSORBNVeo2ow7hVRTXkFPHWa2RK
+3cDpw4hvAniGoSYATactrSVHAx5hOk8fsvQGwUbXTfs9JrcwGn8Muzp5inB0vJm+Ldwxo2O/A87
HRanqTrXK1cmHq8MCUX3x4tJbJnCrdSWzwsckhlHhzOGdIfdcC65hxWjz60oCMuAXXmRhQC9+olh
LO6Bfc+Ii0rHJMuK57kVuKg9bS3ux6s45CWcK6fP3nTDvl15S9/qssgm49V0T3tavtO9FBdhWcOc
aTaIH4PjpOn4o6YTq4pSXY/RSdL8QBjFAZ2eADmoyxo9wUxczpLgEM/setQvZvzTOTiv2rQ6iN9v
VpAlROtTbLRjR3SUUbXFlLYCw6U9PyP7wgfTgyKJxKYq5kai5WIk6CNxzDVXfo0GblXt9XEb7ZPC
izvS5NXLMWhikFdxlP8cgYCoa3Obx9yz8UAnSgjuYr34gFHTEaNnmlv5ZMaI1J6NSEBPi7DxWlvg
t4J3guSYialExJbxS3cgSRdjSXFnqJoRftrRjHAjbzguC8ZdKh1mAmL2hGpS4Wdw7ohSfb2xnI1m
eT5ortBfcMKpvHf54jdwZsstgnC0JLUC4Qo07hLMRbcXu+tUBDUWZ989u9s/bvsRj18cOZAbWZxx
nEaIgCX0z0OsC43bpX0dJUZyzcrOUaGZB6gSON3ENiBX43OumspLDZAtocdynZvmjra3l4Zjxfg8
DPtRvXcM8aKytuDTTNGSCNvxbP8IZS35dSjIeXnSUcp/cai2cjkVcOx/rsTECeNLESXvsQb5cK50
dWokdKhgyLEno+/+HgKevsaMBusMVxbP//U+Cqu32j0GGUoFGfARY3U2jdGNmESxhtJjg0gTXn5W
fvpMp2Tvuqgo5jDWdwuscKMXknnSapBhPQPUFkri0wyC3pZqxgU18oZXWbsz66CbZcXSgDy5B3po
+kxv/ipLhMUEGHrV0Pjy2Fo681Io31dMOaGdLarWG+k5e1/9fGdN++OqOBrJ9qLr+kNQCnP0b2AX
fvumvJTWOa4/WOpdgMvF5ClG+IVYyX2+IkjL0rMXOQWwCEKVsRojz4jfrm3DCTys1vMDP70iKzpO
PimpTDmr3lacWagnVDPE3Cd+Lj3PJaTeudm6U10TjQkCAYE3dNbGP32ar3ib1qInRThAf1sFXgdo
5nIHtf76pyRoh0Czm2Mw0Z34dE2WS+44B48UYjyoe7rYOI/bE6GyQyGx39fRuWQfjTpqD2hsa2OZ
7WrEbPdSMEracA+udrvYf59ujDJnOOlpWekzaRUFswiANfvRhwCBdTUELYz7Y06/wivjCqFiq3p6
2N/m+ouCFxg3uP5h4U6eaEdpmtuWR03QJs+CUBpZRl3Zrb+WSepvpIZo/Y1Ub7xfvG107BDNxDzL
+4Llwbvm2mjxvWa0chymDDlsEuye4+WvDvjcl92gIk/UC3MOoQtQWpiHWXvSu2PT2ln+ggoa4AVG
IZ4LH6lo+BEeu9+Jf1Wghi8qpyeSK8a9xqHDJqeSDyvcrm1711MsrY7jWhLAqesbgEbt0Z1f+m0w
4Q30l4aC9I59GXeZXGDGB91i6gF6xEBN12BTDum6K4Ys4twsKpzl6PyY8ckly8oF0uPtrZ3f8prD
SuD9+C5s8IJAExa8C9GklecuOv3/PiKhPd5DBC8us5ANWHA8ink4QU8uyj+YiVEvZTF3x+e+gZL5
PPKnyg1vmiXR51zhZwNx69Unxe4f4+5yTHFOQqctVDPBoH7tOSx0ImiCxTxUVXEtl3Xak3N8SMjB
boYsUv8zmjTM+qv82dK0jfkU029AtaPz+100s4lfdj3VqSilNLMH7Pk042PakVUHyBjERNAgZ9X/
BThSJBQm04wFLObddk0kYXwpbNb28u7H6BRjgLy5KFPJSCctFQHbo1tSvcrcNqhexN0nW5a3I+ln
qgSGSp8roDHSkYFuYMfNg+3g5XNe3vpj2q0vK5TZvD0ucgftgquCxDNc1XgPUkjK5I7nJLrB3sy6
jqn0JmfknynxI0r2n0aalmW79FwJB+jhH9eVO4XHceyEL0gT4vwErQ4l0DLXZ8G5U4E/DjOfX4lg
QHAUHevGMMOF0HLn9aTnZhKaPz0hH9Cd3NzORB2zxtl+/6wypaEVtfnrluWo/VyHNpJV43g+uCol
dSUUOWvzZmOU5XzvBKwywzgQCvlIMxiAiE/ILoNvfCbf+aRAks33+D0otlC8FgcNIKtg8DOPUxP4
VRelek3P2TBfP63Ax/B0f3DZ803P8aPsxPiJTk9hsF9sgVFvfYFhl00GX0DaVpwX810yVlXp6+y2
zjDd9xhZ/tep6F81L7A7uExb+ENClAesj/WHDaapRBo3tUuA2lINYlAnL30H3aiEq/jYyTiSQdDJ
5o7BLplvvAtSGwn8fqDAJ0sQJFvbhkvJSFZ8AXJaNpZI7EPKfJaNKB8Wkr+aSsEFtIzRSb+GiJ7t
udpeaepu9PkDX2mqsDhPSwhQKfJcDSGikUMisuI2tvUixQ+fasQbmJo2QTEPLptcB9ksH+eEcA0i
YTW8d2kmQRqXldW2wQhzW/q6v33NYVyZjKgOoXy+JiC89WjKSBKnnF4gobigGw5B8i5zlMSjFM2y
S744nFmlUv4xb8VFutbv5AOzq8x581jtCbHaDdOFE7/nbOsCRlKFDN7sx6MbntAYT1gpNE9xatIF
crzQwQlKJ/l4Qk8woysxpIzuHNLQ1GNM9lMwHb5abZUmlJVmhlYBlSFxCi7LulcYFy1woG8F5Yp4
v/e1doBicRhg1DgIHNOO+m5/tCVbty9wFthgodQsEAFw8lqbl8aZTTLKxCQ9ghwREZbdB7Gx8FDq
z0dp1s1QXh+0NAG/L/Q4PBcMA8HY+/B8caDMidaAw4YAKViwUmoWTa1kcUQt0fs3yDMMiU2+5Bfz
27N3UMoB/0hZ9ZRatkvFrxCC2J3JhESQoLNY9kgrLuFtnsrcrg2oe+T2p69uxid+jHDlQwF/o/Vz
dSUj3BO7X+eB41yQVEqjkk1/uayrIo7JyMOtYteFL34XSzcCvG+e85xXUW69PAY5SK6sDJzV83nu
8Iy8S9XBxSVyruAzARmhgI3LpdM+MJcn5R7NdGuell/bj6tqhDgNju09se7lrSQC66GPl+8y6fDE
aSlZOwK1CkpStHC+sJwwiVUpl/T+pC8ZfxLzTOM6H8TR9Bc9lK/AV62G4TPQknw1ORGQC73t6N2C
gvygTo00Zl66HVXFBEJZheXcUzl33luYc1P47IOwYYwYOnS5MbhmYACC9GNgo9oITmuEh31EaoyR
3x0t7BVKsmcyj6LiqS0jtjOLC8lr1olY42KVhl2iFdmLWHxi4XJdhnHM1rTko5qxBt6XStVG0Wl+
aCl1EDbdN20rUvT5kGq6QRulpuE1OsJg2y6kEZmN8shZsevcATRlvcL/RHoIV2Y5qIn4jrQDI6fF
Zo103gTVLbxjf79UloD426Di1O1hb64PvLRKFJmDP0jYn9NGlxL6WQzWVk/ZY/nmftu7/De8ut7W
6hb+f7W8UVoA3MsTh5JWnYhC0DyBuXrLzQEc4TvF7x8qhIi0VydrxD0S9M/nRodep0a4hFXw8YbM
9MCbbpv41YLeCs2H+9IQ8Rqcl2JwGi8KqeITNVKFfqM//s2c80Zc5Exj7/qv2QxfgHYmNAjGEswR
ku6AQ3Rsvg6/zdbX5glscNOEJ0XGHchReLtxORWodq9+ecIibQ3A5g2bhJe3M0uIPinocWGU/3vc
RhPrIT1UfIKCsaKo2AxBCsJ0FT6GgwjDXvugktxrT5KpKkmWmBO5j48RwLveyafmh3oIijXTr4cR
QH3Fw+i9sS9gYm/RCgHvOx06ckJMoy3s2kd4N2LRR8qQKzOr/mXv9CYhgvDVMuee3tAE1ss6PlEW
BnsbBHflWVc+a0KSjB2PmzlgZp4vbXXBr0Wy4psT9Q5DhtvAHRtYFS1YQnuO9+T0KF/PxRpLpRUG
eCf67jvHuWx3bVUGd7YLTVt6OF5R5L3nR8+z2eCnsXY/qN4DFj+tZaJPbR6+ScXTSlRpTOewofhu
uDLVR5zPx83J3j/BbixTL7JyeCJ7ZpX7g4MLKPtMArTSHZS78EIaKZWyKpus0RbuwGvAyuIEglt6
PANUnVy2/jdODAsoi7GbQH7MsLSuQaUIlanetcQbqjKA+5gnBxwX21Uzv3X/Hua2kw1RMK6F/BZI
FoladuQNeRAO4OulAUiP7dJLvhB/G1Rr+HFlAr2kpWFSyaF3KZ1J3TgqVVFaZSRi6lJXxwNskisA
SuMuO9c6jy3PVfvNp1KdXe7A+hcPezJVbKmnbjGpA+z31hLel24biakNWIXnGQibCeeXQI2103Fh
lqu1UhweABI5orKGI6WXppZp16qXAqmAW/FM5eM4tBUXX7aRWuHI2I+9ynxvbwWJaCyh41C56Pqk
uL3VXWUveVIpIatYX1alTOLxaZKT/14zf6AipNGwcIdNU0m6O61QUIt8UoeUnlHv+I13NZG1RFto
E9k+yx9FgINfyQZfLM3VpNXkluDzVYSKURzE7/cmN2LGnNZphV8/fZ8WhpOq746aJhHaLbvFsEOD
cfXJdc9GcieNfZnxoyQQvxKRjWfciBRlCvfLfhAhmeNrvAv2LNwnn2Oj3tcWLzU6XrRZHKOYolen
XN5GkHEhaB+dbGDGREX78f89fwjuim3s57n8fK6QQnfK2H8lYKCmESDcU15dAYTAdpPelRbdhEXN
VJ1cHuwCQN1rWG6srfe5OUDpnuht/RDfKeea14RhleL7w+vpbFNNqG7C/GLyxIaEAsz3/3nNnAKb
xfJGcACK8uW3RAZPnMZ5y7rqLFsAmdwfl9bl0soHeigBiAddmBrdIWGHsl0itRgAsgTST1pvgRK2
FgNplr6GoqDJhxjoV76z9u4mc20tWrH0dof7IRY7muhL7t0jdUI6KtqbLygsGqVlFfOm/srHG9Ea
KYx1kAc5LKzLO5rcH7y05dD2kBMqLJohnTmU3ONjNR5on77vQfdw0weziFnApbdfwsn7x864jRiA
Oq3l5rSRVsaZQYhkA/2SmxcKX9OvqqZ+ijo2s8Cpg+5DlmYp8FBf6zybiaZP/qILJ7VsyJi2K+Q/
qsH14UYOyM2qxxercxPv7hg3QZ54ZTblxGNqjmFtzsFWzyrFd2ztzudQtyYOGHih7CDwCFYLu41U
NQQ5PpOVEkL6lBlvIKhxmGT99Ki2417HwMV9FilB8G5PqTtLF3k9P79+2aUgG3Bql5IGAoKd435c
CnlTF0YpoOrFYoWb9VCAFmKU6C/ZL3AAcx4vR5E5g6S+r6D/0t6KzOXSuQgVoV3gTYt38FNun6uS
q7O2sXAkz+tWkBaIF8OQMqliGLOPjfsauGqk5vzv6OLL5Xe44wCOLahin2S6ZEXERzZZky1eQFG/
ywwutIkNHXACiUAyL9PndRImzB0v7W0cl8Bi/YhCLEcjix5hCinDygYLOhKH7Zx1vMX1LkWmWt8Y
hwnQtegcpwISC4+sTvBdk1vhq8ivZT9NMJSUv/0UDqRL2cJXw1g83zGOssd938DrFCW5kZg8BE3i
VoQ1LibCwkNmLMzb6eUHvBGjFWS0bKpnFwtFRC9Qry1RbgvzA5cY/YUEj4WSi9PdmhrneFseciYw
ZD897Vq1wYaKEgttVs7lDJbpr3UO5JQxeXaa/2pvNBh8ZbS0yvOzWahUDPycYHyTfKVbAp3+deDE
Ez5ZZIXCGLTk9kgxkeI3YEwoKb0IJDhKMuO+qRrj/5CxpzngFfwQORRLBcb/QoeDHdKFsklzMIOm
kz+Uyn52SlHdmn7Q+Xbxv5J1nxWOEoKwLp8PlBTzkhtYqcD3kLGBRwyhPtYsr4lgkZrsTjFkz2st
b7fmE9gPRMEReksSG9B6FGJwzZXvEPzlDYWl5IO97WCRhFYqbaPZQh2J9/cT+sxuhpSEA4I+eiT/
k/Z7+cVMp6Ta6fEdhMnXlZOwEQLaL2/OKg1S/4kRuqP/hkbl0NSn3S122VwYhM1qFzHPM0505fBf
CpLiF3u/Zi1JokCsJZ8X85ZXoWV2pnPzyIoYrdXySmVnbbWIjlXD9YQZ0GL0D8C5Uu9eRfDW8v3Z
VP03nS95m0ZF21czVmpMxJWJeqUjbMsQF6uBj0VtP0Gm5lIAOPIIGwzEWy2BjTgvopQyKq1gwmYL
Dbw5uUHhWHTi6uFXbskgVZ3ON3niqVAABvJu8Y742M0TeXxvfGVT0Vmk+S/mstugIMKHoS0EzCXs
3F7YOxRcxjaDkrbeDfxiTco4KEC+TXKqPQnGC44nHgyJ/EIv6WGv7Sg8DPXmHpaiv0cf/G1ltkOo
0aaYi7Mdu6xfHCmRADSrnJYVz5mh4VJGMBz4JGOP7CE8w+pxnx9u8Zcx51ncGJrd0RXuEXF7gRz2
Uz6lOaP06Gvu5qLzHCEF4kiBS66JkMFGnWvbDpKmpCETZBPo1V/fJl++peMt2ymJO6bYM6C4YF3I
71xNnzcpL6lpjU1x85L/GHZU3Oyxvt0zN+lnqQFttygocmd1AZ1b7sW7WKvzV53PpAOV4/g17vaL
K+5yJyX579LWW0k7IyzzV+VZ8As70BDHgiMDAd+MmqzW0AuhDDC7+oH3y6N9IltINMFWS9Pu3SfV
6rI0jSv2g94jl7JJK140OGktypUxmCWf99l3cwMtYXAzD6AM+epx4UUPIU0zOLOQBIq37go/ScG0
RkE+W+S6HMZj0k2JNT/gx7ecZaXN434SxhXbXRWGbh+FFWcK6yqz2KOaQusVZdm8AowpF7wYMLOO
TuJhuj07Pk2leVkP0EdfM6bIiUXvVlL9BvvEkxoJdk1njbc+7doHWp60WISZJdlNCA/sJ+Z/duvr
1/CSmKWLyuhglbO7xPlSJA2M1HDG6un0O5o8ejtT23n5v2Flf9G6N6zNJpI53FyDBig+5zGjfqXp
JEmcUXfRZvufhK7yxTy9wehsp75mN3rfYhcLcHLkk/uN/DYf27HHn49bKAYAGM1BRf4gTAamNK+P
6EHtdr29k9b53MPxhMYw+bCskylvHCd/Z2ySKcg+Pz3yGUG/vKAYy/vX4JN5PTtMSg+qOpuMn1fd
PR42k3Q0/mjzZCdpabfw4ae2u95jrX5x5EBhFK2Wpxc7nP0f1cLtHFNlMy/5abJIoRRsBNeYK+Qi
qTT7lkpx+0kzTC1ZC+j1kspyRe+JAx6qDIdkw4Fww/WXQOnqhvdE4Vhw/Z6K/41lc3KcIqm06k+z
55KIpMLM6Var23pnDMOkxdcmySmSo3ynTEe9AYD/c+TxYPEwfhcXU8FFMJHZMfykaVTxNAjx6EJp
puiFULBIE8gjtzhX9qamUzc7lh8KPahyhPpiP4waAhz1Clpe6FOOOzHG3e1HO1lqWHp9jh2BTMzJ
zEcybiIyIOsKUGiFm+SYXnMjSLpjaw99wNiYWEH42XQE1xcXp+OXHY2Bm7yJ7E0me8GATDneTJYj
DmrM0tTuF0mtpvqe/nmAgV/rq+X9ArpR2u0XE4v0/4UFTh5RbUell2/KxVe5hZteV2iiW/i2NGp5
JB9olgxuRne643WHQ7gqbLZMDII5SYL4tYWjJRbE4HaFuTd0KAs3vbCpFsVAvjmMKxBmJ6Kx/yEY
yZgOmwug6jHXKuDxlHf78ASOVaXLrrC2sVh/hU07XCBFOBveVNdghDxipnoPm1Mt+UwJ3yB7cwQG
PErrB5Br0GcjZuvuxFWT47/2OjQjHvhYkMYCavMiyGnmVbkeTRLYwXl/iaN/GqC77TWbDfGy6sK6
H6BcMofnLh+2TJ38I5XNro77ojwrKH8xEarHaxNEn5VRCHjpHZBJOngesRuOs/KQsOVRs7uj7Kl3
835ZKuNr/1hif1qbB5MZ1aHJ9Kfdfo5mlIj6bZ33AMBY335wTutWkwQBt0ZR50AFW1hGfveaENhw
xABCYpblExzLs81ZS6KnrcMicoqi6DnKYTFRe3NeMiJaKzyAmeY/9rxqv6svJuHRCviA5WRTgFEX
3TtdMYbqeuye3IafBqqzLAoLDhoy9nUhGij7kklE67OrQvpWmSeVuG2FH8762m+xL3YN0BFhmSnb
XvUOwPCl45c4pNskke1MzVVmQ6P7CanuRANpCWGhvJ7OERurf0lB23X4jKKZ64YY4va/pg6L23oL
KwkLRXGkPsomeSqUl2iRGdHXvhZR8duTcJUPjckhruWKNTVxFcXj+hlPC/TabYATNMXtx5QEjICc
NbnOREXCUfCRlmWWPj3m3AgKLG5NfDHlinzGQxLhSAMvTTxMiCA5OsUI72GDcM8ze/jU1XXY92qk
b8k3YiAnTJVFfpnfsIOwIaxowqiz/k5/vVAgKGldNNCyBrozcyCjMQbS/P6ADv4+jjG46sd1WAUO
p0r2/TtFdM5XVSM7gfwgzkLlNc5TpyDN1FRMoGxLWMhFwiOiBNFLvqRDLK0TQnCyNkd3pmYWsV/C
iIJHvsVGlB6y8oYYGEUDrDlQAtCHJOeK2z4NGGPEyvXWYh8PAxJD9kqSdz3x07SI+OfpeYrbwRsI
rwmB52+wHsFQfNpzRVNldbmAYKl91KetERoILPU79aiprt5rRAPQqvxDESEPwMmv3HeFtGLQ4gNK
a7EjJHhcdo8SPyAavclNjPv9sSJ3ovNlknuBUDmhVsRCQ+02HXdWhKtvAeff6ahSAbCsnyW+cmms
XpQUjj390hq1dG68fzVv3mZaS08Ndqx/oCjt8uItu54x4Zs8Ycb2SQwYghLBPkEx2+dCA42VNvei
nVgpP3wu9Sp1WytR/qCJfaUyJI1bbx+m6iD0Y9320J8kaYmkoaPiqCXFTe1ikK5RVmZ+lp4y8j+0
Hn6g/MbGXdVA9dKLKpY8zj5e7tkqW7Mcds7LoQLR8CNc4gew5zH7L5qubgkezCNEdymf1nSJLKiE
TifPgafBhK5Xq5eKycrwaaRrL6Tt1vEbIIy+2WpEaWXdfNQ27smKeZV1kNO8MvJi3B4T5fw6LaTe
qRJq7ULAFg5/S7njH3KQVDS1RHX8Ci85GGofv4rQr79nU6bfkKLu13xD/vVe3LRfgiEYyEJrlx6y
GocklpNVgLEMOiL7tZXB7RqYFbn+9zhs9VwSl7teDx0i/i6FMdvk2el2LWTw8joqNngrMFIOY7N7
ztZpaQEI1dTbkTJo3/sWJgbIV6YhG3QVle1plBENUmVfSxHI9t42pr5qmY2BqcFn2KK03kBayYPf
ylYD2PeEnpvM9zmPQ3A69SLM0KhLanrTiL2SSVgznKLIH4tjSU+VfuR2cv82Rb1c7bf871tg9YhG
v7GALefY4YLvXcD5UdXr8Ru+HwlQgJXrDgi/i1ZIHhrLS6KksQyIq3Bvc7tJpdaSae+M/w0jzxph
/VDAOm/r+lQnUrCqMs3Wh+srBT+f3Hf+fNGyNtzMyyGfz74f/Pq5melNbnFRVwjGAqouWlZNAVL/
lNsZDZJPfn/oPVtGVoSrFm89B97o9YIH6l+Wi/psB902qbnk14oryFw9UOPu01HseZswPE4tq82h
osv1G6u5v1uwX4F//r85eRyO/OIA+pjhMH2FNcNH9jMucy5OJXAgCG6kcfHXOj2i2L4JkAcTn8B9
itLst0A8/zVPgvUrnZmTdQMZIqDTAeQQ6poguBOenqnUR9IqvnVi3VtjVHwagDx1FalZgkLUDvmL
2+xyVcODxXr8MBDpz2ytvijmZKCUegR/s9LmZvxinsuJUicOARL6OdGv/5ONERJxBbE+cloaR8Ob
CzX2wxKsFcBrN5MPifqTn1tlHI/GZI9zKNCvnuGjh5scD4x+Ivj1Himy++fYq4xgJuCQs6R5+bAh
snJF2CgmtFY/Q88+5tMUWtRYrb4VuTxysAyd/KpxErhdrhZzHdAyHlMOvkHpvhTeyb4JYVg3sqWH
JiUyo4a4aIxzEd5dBSb3VzJTF7k1lfmR/M4eFzbvQJbm7YM+chI18atfZReLnHaQnoNDOaUYHrU5
erxrxfcAC9EtUVL2jImtL0FyKVkT2WcT98hQUSdY69Eu/zBFleeSRm/sXve+Nzx30U9AqRl6eLGp
IzsSyctIaTQ4f0fS1c0Cgdpq50UOr//7tNOBUBzeJAxmQAAWTh4ZJzuZwa3tbeIoZpHQoHlRAENv
OG++XYuPZa8hZVV3Ys0ZVwUuoVj/o8JWnPrPFOpns8R0PPm0qQszNAENy4K9gOU0arxAVV9dvJ3z
nCAutoH5CX5pBfmtVMdbPTtHC2xM/VZofewlxiZQKjV5Ly3CHR8L7Etl23dgGFZtO+c8F1+eAeMU
1J4AXqEn8VaDVMTPl1uiY2yErfxeM2AUUWCjUhdEZX8zPpBIofH4tYGU3YHzxIn/V6E0rEyu6EBj
211RBjiSZdsRvdLfaaCcdcKUN8oqPIPWEGrU8tdsFx5duC9Q/ONKul9pmbMnL7stmWYE/40BL/WG
A3JOAEE0hs6pobMo3g3t78vdAkb+aona+pi3UJoIWwJQr5zsJQSVy7selRAtFe1Tc88Nkl4ggKr/
uu8TsSDl1N5qyC59dnQuTPakOpxPFmzyHheCeb3sslPd2v4cb0WdlAgtE3bw4tIqxo4mMjUujVy+
3h+9pekh7yQQpRb6eiOHqnkKYJMrBF/hR4iiFw728k8xF5Xq2iJzziiPTd2f4nlABdemsEhCZMZj
d8l9MTFZNa+FeCmyvEloeiCLnE13KU1gU3T0tjDBTZc+QS2H2Y7zILMQHn1GSIKQYo6HrGeAedMK
u8q9/xhujG/C6wzPHb4cCf8+9ZiEeFE7g6/D+i6KO06pHV5X/VoXO9AXTvGf+xD3T2+XrVwCFhAj
GWpvQ0ejAaKZlqXSS4EwNjixeGxFJ6MehAp7BNHhlzHL47xHwgI78f/LPhasmTAvAbxkKdgorsGo
jWTjkCNq12s203NG6aopo3/1sIDN76tuYmwy+xzhYb7COwRw4TI6UBNeUJVxQYeYlNt46D7nlVFs
NNJjEk306Jxdk37CytszrycUz6QORiJB12KDmyTNwzsTamiV8oGQ4QhSpBGb31cK9RZHmsNqdvlj
ida+PbssQ8bHw7JWU2NjI64G2pyiPuLYvI0k/dMnEjVcd54XyaaCFbulxcww2flhXsaoeWVVL0YV
3GPHVNPgjdYwKzQjOlqNSLxIxFDeymnQLkC5H4C4aUcKZfsj1kz5LTjwoDjVhb8BWCzCDXGRZ/Wc
i8rM6F3EKG/BX+teCVB0TazcZA9k3k0986XfTZpRGChqppJWn/e2G4p0heWxPD6Uyli3GqopP57o
Jl7UbEv6VZrNHevsQpOyMzM/YckE7cx7b/zc2jcqMYDWsTps1hxP2Y2SSTKVPOx76DlXyB/f+LIu
Pt4xcU+ow2mqEGh8yEpuhwBBu8cZaPD0ZOgazsC3ZP+36l0Nr/MCmRIXa00U5SzTMtzsioaZFl3/
J+x9Kp0tTveYkvkySIU8/RVYu+xNiLWkLxFzQ9BV5sEi78jBEK5KGsPQ4+4Kua4T/UQaojNM8UIh
04WjrNQyek0dXokkOT5r1dAp4YU5YHmyxreJzSH2lua/KYQGwWd8fJJCYuFzpPeI9uI8Hve1AAJ0
8LNPm1Fbb3CYPefA/pcj4FY4PiuqlaYUljjLGDWl3+ssM0X3jkcQjRl3YhBR9BM2lOVjTC2dm5v1
sHG1T+iQ+VjU01ogzX64JfrJCWLceeHek33bgjGnG7b9t2ZV0peOrg40tKggpR78RbTSoZh0hawv
QMh8Fkksnw/2UflhQK6dN9ru7QBXp/L5TOhVs5flcYSfcZBbNi4wf8KUerik0/+eR3iDkSXBzRoA
/UCvAuoBy3TAbgwhUzN1GQkQQYimkYEyAm7w0npPNBevL+Sb0TaeEqRlCqYatE3ehKYnWWzCTcVw
gvIIAP7542MvDi8f3uWMgufjrUszNFRzzUImXmyyl3aX+aXN7PeIHF+xMgWuJouffvisllNaDX6V
Y57BIhBnWcu1Si5KUPIkax+UJV72cP4N3AmjL6X+MSIjngEYIvxi6DCR+WYeiYF12FcDZMl/lmOY
rQhYP4asSiDoYOYhGvkpT2deVIcXGuETN8VDqDp7UQirIlmY6Sp6+x+BwcTZh/rFT0sIDLHBmmi4
V0B/5JTPQdFasZ+vIOMp4YZAhuSK9I+ZBEwnTEwjbH+C+yl4FUijHFQjbIDExDBTZvD3KQ7X7C1e
FC3uw9TqH3ThHFIMf32PAsYPr1IU2GmTXNMvqriYPI099+xEMfqQG1CngM2/8FvWDrd9vyYGfANv
IfoEJHYrc57Rz8vbrzwcqP6N1guaBPTvGbLSdB3uYjj28zz70oAsEsKin5oxvqTHFa7ThoHlNCxy
8yEie9VTyzCbI/hpRYO62VQQ3DgbmUxkZLrsk+lPpFG5DUhsT9h1AlsUgYDdIsnw1w+dKLdrZ4Em
mF0cSS9zQ5ZjCXi+KGFG+e33UNiwJbJ1WFTNCu9GxQbARlcmAQsyQI2XgdSj28+6FP0AtFBItAsE
/CmqcSnsgQM/rvk3e3OO8yBfBPww5WwYjH1Q7fVWWsjO7NzXKQeKSFJmFb8GP7hNgoC/8iY9ysSS
3G+Xe1DGV0St24v2MVD5iD4bctjpFpqxMCJLEg2c11S2qkeXQY01VcdqZ0t/4wsvdblC9SXwJRyH
X8GGfQsoAOKrkZjw8NR4CWFm2fx7IHDmmpu4ev3eTG6EHbwYH40xLspY3ZagM4AegLgw7VfCF4a+
5xbutqA2MWi7pMqravK9hB96RNP6xfDlnL2HuYp9WgeyvfoctF7Al2zLT0aPNArB6yHv6Czw/hyT
D2XsC/CjM9bbyHH7X1tH8vLEl4pcgQb5jLxWBECCs5MH39X0o+L/4UEiPoxxGZDc8Q4VpPoSZckt
S1xcHwUJ9bjJ1HyPSPB7tMCZGP0toaQfCKLkSfRw2kltmVJTm3EsSchEMUHGnv08HUlWe6K04Hrx
U5a2rgoh3o50Kv5fBIasoJo+LPBg6EcvBcNb8h8WWbEK/94hmEI7UdD5P5SMy9j58pXi4NZA9NMk
cBycyvVwsRoyvjK3kUJFGw7IgW8nIBBBP4aF87IZcwQ58jsIqeYKZW2Hieq/ENOWzQnMKP75D20c
eWv+IpvWgkg4orMVJ0vd5cWztsp/AagL0EM9r4/LkJyuciA055QyO1ZweLzp22KRuYKNAoaA2dox
iy6nAQ/7O51/Nb2AigfUHaKMke2x6hEWsAFRYmKcI3GR1Btyp4vcvFxoMOJWy3N7Ga74P2uWeJFj
BuHxGSKeDSdkBjzHvc5720B966qOGwG6KvM5KKqsOEPqwOOuY9lUvtljqF8e2CILSVzPeoukQi50
WqWfOhyYVR0nHJKLj5xJUGDAODPo4yu1YjzgMsmvHNzzsiNRkdHf5LgRT3Py7z767O0cuB79nT/j
toHZ8bRRv7sTsrkddzPBxN5ca/RaVefQhvrCDXI8DNEU+3pXQ8Cy7Z+QHtnmonkx17TSTU4n4ogI
+cH+R6FONMZsX8Nbr9rx6voXFwf0cBgewHVIBdTKdZnazZTZHFjBF3M8DC4xnFZnD3zRBC5k24E7
zGuiNSTS3VYxNp8wf3M7/NtWTuCygRbLVkA8TNFMEjq2yDVIX6rghT45a9cZtqa1LyC4td1yJ3Nx
g6NQk+0sk3h7oXOkk0lzyVhR1Kfb82/gA/3bnsqoTAD9TuvrOizEjlmhzlDCMEyez22eAY+y+quu
ic2QvGd4ELlxw1S0N97IYfd/KUuanvB/xh5XcaM1sFolblH5BdlS8219BXqRxsstFaDGQRWH136T
WT+4zBIV3+rXYB3V/Cr1Yo0OiwDzcZKB1JV1j5rKpAdhnbc7sZdAJRNgiOWuoQYL+06duM1/YaHM
n6DW4cRorf69/FTfi8vSvXLMRvvlq9zqU6b/mNhrYbp06Uw0hU4ZplE9lAuXuX+CgaCv1eh9dZ25
7tSQ6Tfv2MNwetQKQQyE/cvJjsVbBcVHDOznmAmKiwmadqBteMPILhcbIWmb8eH2vw5ePZmuf6mh
HGu+AKTAfzSqrI/H5XxoZfK+vDxfhIBVq0rfTBcmxlYQn+BefavJ2UzgSZRD5GaWDEsMdqJdPsAA
0f8CP5igTOR8KkVPmHlfLedF6tOxcbC9UglNS2Wuo1PtwBiKUo0E+CnfmhFAFpFv4UJy3+C7FYcC
k3XkaeIiBmFx5EAry91CbXQk/8dachFtkDMsqMWPt/FmpDeyvVzujaA8JHLnOu4/57NPJvzEwYs6
KN9NZ6tsCur6lDiagTAON5RvLMgzM7lejpKPZhefpjLwMzY2S/1vr2n4OMN1tLzDt8ZPf1jzRvqa
8LXelOFvS6R6ec00ymU18cjc1naiXI7WyXSdKpepJJFOC3jYPL6GzK+k6S+vpaLq2DKvduHyjXeP
5rmN/Yl/63oUJoEzqLvqK0ikyM8q2Ai2qHmWNYexVoebU9bYMJeMtf4I8NwDH+u2jlLqObDcLbhf
1l/FhFF+uXxe8OslJCz8U8G0LGhIWJFPTowBFKu1nt3EcxapJTJgwELGxdNtYC6sFMjMLtbElnnr
ofgA3mXCNAQwebalIeWLAQReeZD0BExONwX/3cgMk4fTzGwKGKVlvON+wcPYeg+Ka/AbtVWd5Id1
uBWlz5n+2mz39h/TZrtVtf68s5aVJr8Gxqz5G2rSRuVMU88dEfyFxVqbJtwdhbx1nYzZrqPWCTnU
mbNxlSbrmiMjxvfMpjRg9bMNRTXrAsxQiDU3rMvmXnbfG6S68D7klowniblFsE5QZtY9J0789lup
NSjw72zuGP/kWG/Bbt4GOVj4/gp4Yduzfp5QMLCilEYssc0Ka8VBHBJNat+z2j0lPuxTxAobHT3y
L+tn0ZNzu0FGm9zIROMPwNVH0B/+1g4t+leZyX8qe2VhwWm3KFobJKwlB1jEnNw2hGGvduYKqDlL
QwbZRhlT2cq4QX0ZFS2qPIHe4lOEBCcnclKK8MdTBnawICpZ6Ys0KFqP5p/DljOg8dKWDa2Ycwec
tebG2sfsuwREj16n+I4erMD7OBiDz5wrGeYw3InUVB3K++VTvaFUwcZtvl5mQDFSOQw8IY9Aop7f
LTQyNAghQjTmI1n9wwmr2FDNn9wsLBYO38tQDJloa7kLVl/hBUgBPr+A+zzWMMcxNvN2mFbhjWn6
OAE0sPYjTWvkoGUfrX/ZuBvjsdls+lDg1KCzhmKvV1wE2rQGbvk+YT3wU+bRP8RJBqS5eJcF1LUO
WFrnMe2K3XPHOxcW7FqOmlCosibpdHMOShY/yZKie/tgcZpFerjGv025sZQWLgOHYiWbxO/hbnhp
gRHwZT0ZM63f/pJnU13jpe37EWfTw+YmRHsw8J6/5D0munI1jHnZeyHjdnWKiua+7f/qpZTJHl2J
lczIUE9WxawNHfHfYDRiN4zdfW36MHpEqj/4+46YMthjN0k+l/TlfAm6nr7/VAKyf2xi0PVzrKCu
n7DwGdffU7LFt5OsBoEmQ2+R+Z/nLk4vSYChJX+wh8fMftFawT5pof/sMOoWFL1JcwXIxv0k8Mw/
ILck4T4LaRKuO/pzGqXwSg5JlldojI/WWFSECeEow93b/SuFXI9J6YMHQnjiKfkV/CGlQ6CDhbMZ
zPyAfFPoaBmgb15TSiTnoB0qbKyFWpSvqxj+46yP0C/3W6ZWpUS3+vHKrL2vpDXtLzwDU1CQScwR
taPe8is4LtsUXpORl4wTEP95ZI4NlZZIF55IebIrwOh6U/61YJxenDEOLuziLNKtYx1gTQvilKr0
9GECqHFOPPCH8JqVAA7d3qr0pAMavsyrLtQnKkyzd4DTBZvHfdH05E3YTcVxi+92R0Myt5wnALYW
PsbTZNZsHYK2RFVuz2uP369ZKmZ5JRMAdDnjjW7EsQojSFmuGZvLywoXNG72g/hH+hnnxN1Ij82E
GtybDpXsBxKU53s7NysS6VrrCLWXtTCQRfE27LmEtiJatuBHLlo/6Mva8pAcDqL2fgab34Dyl30r
UsszqawUI2p5g4i97PkyzqUOnIXy60UhHQHVAlqW5+x83zCrorMjUYYiaq/WUkbl7cT9TN6VZ5Cn
NjrCb02QONX+lxCzFrYyO0k380hG51Ksw1WtELljskHDa6nrOg/58p+Zaazxu2mPiLBpKk4YwgG/
uSuyKal62CwXxqEQpAAN4n+x2U8nhaSUBjI54jxxgj5k+qSEdpRs2fVhtS46lPiXafqQPgJHao24
DE+usv7bkHV/QI6zJztedDLYf90gnmLl7d9OarVW2ala0rhR14Tt3x4rF1WpHrgtG4Omgerp45gO
3cegi6I6oBvGPI+5DPPlw15V6ZacZs6RG412CHTL+MeShFlWQ0KvGabcqVUqttsZhYogxtjGCiJk
60eVqIwZL0Xp2VGKAlJvxJSsf6ztuNsOxg1qsLXr7j8aiy1fNWkgS2ZksHWcDYuG+Vr9IAOKq9Ja
VYvRSXNXbqgxj1f0s8M8VZtwFfQxRa4oxYgtRFbwsjy+4HIUX5uk5ML5JfaLJhNWCQ0dhgy8HeRc
nJ3mIdXAro85SK6ctB3FzcBnAj/kR1XHD+IuKUQMFlfwsALDQr0L7lvvthlKGI8/jm+fxPxqgXFA
3Om43wJNutF1yJtPfc94OMxIxBC4U9qBOo5B1eZSdL+g/txMQ51N7S388DS3jaT1GILdrcV1Y2DK
A2A9Y6SX47r36QDhOPFxoz5CUwo41e9kGmCVEKb7qp5oI+bZva22G4S3h4pmMB8l4lTswhw+nM5k
ENyb+PJxr+V3l1Nx/QRinbRGz2BXMJ4QTlFz3jOuohKk8qA80bBInyRZniak87bbnRWL7eKp3a/a
bc1HumJurlDesbq2LeXIGWmtbnsBReMhCTfEfGdeKdaBCeJF/iL9td6Q0gTnhuc8/t8WUbPGq6SB
0h3V6JJlWYJEv8qiLgGAK2AkfQ/0HA62EGUoG+GpS3TVXHbAA8DlVEB/HEehVD5jo/gB3jdBUi7f
ePw1YUiH71+1Wanfyp6VzmyJx2pSSo2J+gSUMeFCbeOWEhbfScKaxPV6bq1cIAu5G4zLX086whhy
WNLzbFZYgdoJokkSP1KGfFv0nLELaBB4RUQwRurKmSUy7zFvZgKDjBj6257aADMPJhr4irNLpnOM
lF9DQuVvMs7HMnmQI/EyjBUo7/Rc0zQCPCfz3cPhsGf1nrJw3acGJWxWzyI7yF9B2xTtXk+uQoHE
WW6RfWWTFszUAoZflE9hUIvsZRBX5pZAuMQVip7zKrqtLCLq1d7DS8CVCfftHeJcrSagqcTutGcR
Jf4AI2rNxObGp6q42hUM4En7yj5ta6BJgMfVEEEN/rbtqvQUF/9I/24CE0E4xFkBGkXRQ3W6WZ2K
x5YYcsDJ3+rQUPhRPE3ucGEgh08eKv7ZbXb588jL75zPDInThwhu0o1aSNMH04yvWuCu8gQBiFW0
yJKgL0TI4j7+4+40ELvoWPZkzJJnQDyvaPWXtPaXXF/bFb3XEforpXRpRl0IAgAbkN8HoSsR3yue
lytKoTBEy3zCJL71aC8eYTYgAkKofGRsNE3EOx9VJ1889rdlpZjdsyw5UUb2B+LPSyWm75TqHFjf
Mb3BwZxCFZBgZ/bYHnpV/AovIJlWB6IKJryFjSEHXRmWW9KrHDhrgs5JAv+lQ2XB/BOSLfAK6Cfn
eaMNs2344l+Ib2EUj9fp549BC2SKdzgj6TvlEWRe9SREUYI6NssFvolRKAPvHCdYGShSt0CLWMne
kH0cr3omRo1CMQ58HrZBTsPD71WihUXTHta/VtdlwIXtDSc1iH6B/iu1iiNswgY+iOgT+hWDVqLB
9hDhe9y5Q43VwXjNvlI4jyXM1zst0lUNfAtK7TS5C9uAc3WYbq8LCc511pkczgVEr0MUnR0hBuF7
x29kFtPF9AE88opPT5L76g2Ph+YsfiOi2IwiKMkPsaI6wuB9kz8XB9n2oCocp0kKvB4Bmh1fEN2y
dTm7tyfBXDyz6JzO4FO3W7gH830auXiY/Zp2E6Zm9TPNTdTMAsMJfUahCAiphQekJw1m/aVGBrus
14hkdy6PpQsem/xv7wPmwvWHiaUjt11A/Z9CtrLcd/drfuEj//VYDxsBSdaxZs4k3MMAtuuNksHU
DnXAVb+5l8cF7WOAByQLZccu+IbvJ1EyC6VIjW2Ck5vTuJRhs4oEkgDhd1PxHrqzzCKzI4tEfIQU
WFJ7SCnuTFJYbMua8s88yYwb9nFcFFHdeNKg+ebJ1YZjghv+a9r3zejj2In4xOa4c0470vDl0W3y
uaRPhY2UuhhDeCaPwfe13RTNPBGu8htv+7WMfxIArP8pcZp1NnBWiridxBneF+2tSyDVsZNFaMsf
Xp2zjz/H65KNIZHBuUsNtm9pJvKUo57xTGdqIFBjj4O2Bxo5XrLsDG5gs/HXwd1oDFN80GrLvGvP
JmAxIvreUJKCPCdHb19GtWEy7vm8nItDV2B/ZhHWNj52l09MPNYQxB41hhggT5XOR+24tMMax3No
ytmQBSw54JvwhYg9BC2373vG6hpXNuVeO5681CrfXyXGjNu397WYGZL4szaJ5sCTC5iza86U7own
vhfLDLCIs3lI4gwzpxcYVZ1n4kCoiSv+tWAaDgB9ySu+Rm4iJ7xpgl9ZBru5AXUasWeyVAxqsVyd
1ONE+bixKcVzRwtvL0gpKMr3ZAwvRHmaWCR1jO1so0VFbBlXbkBkIFE5wGbCKNsjXK6eW10vLFRH
vSHWOdJFkK4r2Jd6q8E6bF64gjj+g81RgW8bRnAVy5V1hw4h/uOuWK+AvWyD4cfmd6rNUsd4vP2k
JxovcABH5vU8t38g3eYNu9rJLN2e+kBmcOLV65RGJRKCs8/CdO3VhnMoQL3L8EJfOOzPkLGB1dWL
ka+o8Jp6UC8ZqeBwqKK8DtjJJDTFILSbMXnoA6Wp/RfHYLMf/tTnGbBwRZj+4jRpI5lNEeUFxgVS
B/1feGoAQtRmCuNpQfurEKyiJJbPj3+VhcRlS5OR9H5GStnhO5BEOhZVWY53CQ8GOjZMSAkdLNe8
zhMF0mPr54092U+Xk3XY8PbwpT2MGJsItZHzH0FFgDeYcWHUoYpEc+rKL1rHJz8uU8P1Kvz2T3kO
UaU5vewTJV4FAisdNu+tFqHKXSVNWAP4LRalkGAPbhuLT+aOLI9MbpamdwKH5q/KDMAa7gOCvJyc
+ki0BSsLOLJYFaxt4GQVX3Q9/QlMbIC1DHdqy6gvvVaTWop41zY5OhUHpj58o+Xp85RVlwvv189V
BbdZ2rq544ewzerRlW8kNDh8cGcPif0/1aHCq2l6rmxnW6UskJpQqE0QdtTm9/E7cTbZib0AY9gi
hIZJqCURolwZGDHsouFHWiS+TNrtV2/WFlqiA0emot7D10IC8uO1ddjXF3+gccmu94nw54ouSl72
FhErZBjqak8fSU28fxzmP1TQH9bP8E6mzLFTCMXFWoUU2QUIy0Q8zX6URhFKGGObW/q8+mBpW7Ei
MJH2zo2FZ9xWbSQU5yy2pqMGO/FTUFxjWcUIEl10L29Fw843a9mzHA0qPwkwQRbPYKSt8RkbQWGP
0WmrOq/Fzu1XfyU01+bNyGe/3R8U9TCYyCj02L4HlEGlbzOMFJ3/SAi2Az/BWbTmo2ASXks2H6Qi
PFehhOMaJoQ8GOM84UTEaztthn/9/dzcNbr+a5XE6UmjgyUbd7EI178YqC41Bo+Zo0f85csOik2y
mKat+7+iQeFdW3Oo/AKUkyXd3+NPSadOK0bi4XTV5VN8TgPHNDWX8nNeZwmFGHlgdmbGtpYNOURp
Sdy2J+pJlYM7NNSe6i6hkD9yLhrNQIZVyBcolGXuD11ZP6gBgUX0r5+MVjVxH+lCKREu06C5xgrs
1f6DKktWHu2MPjTDDY0uh/9L+aDsr0e4XkGiM7dq4cr61L/MoYdexQlWSYadyA/AL9VOfXL+4PNB
AqZ4TKlwqZqbb98H2/syCgMBEVE/Gv1j9R2JBCKX8tnD9zqSBLawYfblY1NfjGj6gfymnfDxBs8g
10GJp1dbr0hDOWqlIFYRo38tL0mEU+eMy2HYRLwi7RkDRiJTkX5sMOFux60SYivrhF3Va/nE3Qa6
UNt+yur/PMO8YSpI+SBWkJ2nakgM3uZAKlVQSoGVjVoTczfAHak19hjqQuRowt+LsFLH/PmhG5iO
oBoLRw0lG2oOy46nuBafDyha5C+R/m4v+UfYhDwztveSHeDSCgcTncdageAkbaF60gKJJ0uFBN6f
zoxThRlMXRA2gReatynvmlpO2b1qMMXvSrmmXH3HS7+L6KiZimzCpZAm6490vM9W80Abn9jMggNo
mGbRVjb0YBpgjk0LFtpSNqUp7CnIC7cNNbw2KxKs2RyithIJkvbs3O5VOVgyd1kRsNPMrafSr4Z2
Ce5AlUryH47O6tMWmrZoT5R7gYs37bJp7OH9MKPfh2LYiZcePybsi1eAyb2foPQLxHE4/6/HQ11C
W3p35/a2arjUlnRMAlC25bbJgZpzTLl490TEqHhtZssr2NCs5G63aD5dPEXEXZzqQr0WJRj/87AO
DuYMXP6nKyfOigrP8DGebOx8VUvcfqTMcPS520wRo8GXCmUgzwIVrEfl/lU7bLlvSPejoyJPzosT
BbKi59hlE5iy7pIq8HJ/PgiVMzIjxzodgLgpsUw4+jxDJyxBdY0YtjpSLuyGI/b5Fpsi6EiZwze1
uE023hWz/tIdaRCQeHAsewzuQZL5wiJBi+OuyOFeA3C9dO+JD5jjV4iN411pbSYLTn31as0DyGHa
RX6wp13FUxM8CRjbxaU6iLO3tK/QS9MR6mAj8a0H9rMWPRjtgboUPAUyPporNS5Vw+H54H8h8k7U
2v60tdUp4PWqk4xKu8E7OCeBfqdC3ya09JBlf3G+5d9+8rY3eABj4+ZZopwaNm+lfyulZL5fCPRW
x+JtFdsFzG3qxE0Jj0IXBiVnzqb2YubfMoVJDHeu61L2vWqUUSZK+JzNmjBT5wr83P4iDh5+r/qk
ZX3hdf2bPBUpBhorlTUFpC7WrvTMeUnVW3xbSuIyjyUr7dyq/ShBYRzzLSIDRD0WHSKC+NGWR0RR
uEX6B7o2UoECtqUmBFLMxWlIdxg6sWNx/eOmoh7yWa7XurFOUMS8s7+ZdjNv5+Z8ftQHU9JTJ65Z
ZQIMrkZYhy761faE/KzcGs4w1UXUH/CtUM4WhGRVRnW5SXjw31bX3OHAUNsg23dsQ2ptv6QYjnr1
1Xp1DmwjVo8fgUQ+E0QHV1cqSqd15TeoP7/P992Fwo2CqZp42Q2GyiUm5NS84ws3HbXAUkqHqGdx
mZ8/Ml+w2WRPlhIcoIKGXHfSjfm0uBcbtHeua07zproOxU+MzNSpoQAvH58TuEaPtqJVyIYjHJ3p
Q1tv/7frJTR63B8Dey5+mMMvdDYZBY0gbBftOrFEoGo7uW6wceQJ0wP5B9eFrSuyBc7Cg5Y/BIzM
/hRdnax3dDcT2ezVr1STfZWYQ8yeVBWgLGALV9F5Avi4pPR0BBSdGnX+cTfglujkiLLhc0LCKaSY
pzDIjlbEj2VL6Pekw0lqUvHwYvZGCmxxdqPbCRrytYhYKXzYbsBcCqRR71hmJCa+uMJjelfI3+Sh
oL5ypHk6P1lWAznLL3tpypJ5FsBNqb8KEQP3uQkeUNiPzdSfGI5eAfe1Oa7DhXe2tuVgAUxVJhfJ
33jUGz9uod0CZ3LF3thtb4p9v19rQg+suACJYhYRm/r1d0iyjom8jWMgODNQKzt9QF5/jVi+yKge
JOuJJzAUwZluuNXE9XWAOTebWFEm8JOGa1YxjkX1CW7lqUfa4rl58qau9G0/SgbwvKOfT/urgi9p
lGT+lELXr5iVJz33dWjnMkqZPMzmPN6vQolpF/wUqA09X1nnwlhl8vGMcZEyX+YTC1y4jBciXfZ5
SmBIKE8GR4gDkSbRilj/GDXdppZGTsg9PMIkBGR7iyd3El2f7xTBv8GLQW2cEVTMV0RcDam8wfTL
CAw5/5XaqFl5awLLbYLa8DgRbYnVJZU6N2xx6GZOzBp6nMvpBOSwVz3PhNplZn4PYkijIoL5fbzB
HggBSXE4peLI6dcHMrJ+8tBhPEhF15pAKWGOrYViXZkvgFvkC0GZFJvEUO6EFPPbVzkGb7nvj9Xb
VgG4CLyNJzHoZcZy4s4bruQ2fjlbxsyHeFMrOnUh7GmZWTiY6cAHepcCvOxiT15eDPR1AmTxx2Gv
+Srsok+M+0oXIzOj5pIwN0OoVwIHXwNeMw/88xzbkk7KIro8c2O/+bgLOWKMFsEQ6VKNCWhL2WnD
c9+7RH9WApx0A+0r9NA6+et3qnZofKzd6ypiWhZN/dX62ZKAw4ZfgJZaWN19BqaXHyCk/WpYQR36
tB+ZJJ6ME9cPwU4oQI1m+uyyzcc3COdRev9D24zMt4rEytFBrpngZbp/6OvP3nx7TvUHEvG86gCF
AcBGJIgeGd7whhJ52FAgQxK695N1OgzFCwbKujVjqdTSj+NnsHxOBljcl3snSDmM9wB/XhAOohUo
b4nXChunFTRs96FCMMFR6KnCYXiDiLJ/4UrRHYDUWIYKoKIlIzBvsF2mDgeUlYiEkeN5OFwluiAJ
qnI41ZoZ1xuPdSUswYppMyRD3plP072IFYFajNH5DNitiCb7BU1biwBtUW+3jmejZ9+JjdTE188s
USc6vi/ELjbipBhfcofCoDDQKYnOLyI+pVEIZvpEGWPkS3Y2eJ2OHgEBmifJ7OM4e8TXJnpjofoX
g3HSIhl0pgww0eb7jHzwUJPSh876u5hN2q2f6E3f4YejwMfbXP2t1bNqmJ1iuWMUPedtkJT6PMZu
emboZH6XxOR6s+tFTeN18y+JDp5DDYuHkZ7f3n/zBPR+2J89gouqUyGTuZul5nu6lViro9o7awx7
/zGvwhLOl17Ljp2VRPOVvljW/QuJi6LOyI9Xah4ZIsom35gGG9iFozFjCdfjEN0kOPM/LFK15qZZ
OQjS+KfpfnWsS8XoBFO2h8xRmeTQD/qK8w/h3oFO4GbkI3/GD2AejsvkoXqHPULx1OuJiyKR1A60
N0SV1zv1oNLQkvCNiXtS/kTtmcONKLyjCHlIfqBb1i510J+Elf0+woXfNyHqIWWa4lltbcDgVRE5
+cemyvCGOCw9Aj3oumxnl32uwSpGzg5/8jnWKtZb7wB5K3c3FtDeaVVHvDlS2Sx20ygCHNctCwT0
7s2687BuHFfVMgXNDOmyGqXFHU2ns3mqWaeGlzh/yuhiwnyw9GmJjZOIbdeIAi5B6YC4bHx345Qv
Laq22xIzFzZq8G6AYqP4r/iaEIPm0GNudbfKEr6DvoxC2sJMDF41AU2rUAnhvgWsXlVN5vgL7TYC
MWw2O18ASDWp2GfUe45bspFy7mUPmBBPloIpKek8AS15fndWbvUIOjqTbci0EX6xJmaUx7phpK2Q
S9nFBq1JK+b9tDQDdqUog7btr2K4NQlWuvKOlfzifcScK8X3vc03bl8qeL2VbJXpE10VSuOP0hb7
eheodwAUvV32fBtN9Khw0s/6kRxP1pu7EOQyQOD9rVvh3RIfUZrA/ZN/c9STq3F43npfwZhCdEfU
rF2n1SrbAZnIwy5WL1vjrGmUU3uJVMgALVxtm0iARBODlAzeWTv5sYUeZ4Ys+K3xabRZ/2aOhEbB
N427fypP4KfjMP1D4wWuKIXzN6J5tPe2LDVvphHxcWfGlGZhl+kR7mNeUhU4/qAFCe+l8tCSbfy3
rD7mdYjlrRGnrI6bkLwZoHoumwMnBt1Td5rt4xSvuhhdw3z3uDdEpcc15AiHuEsJIne5VIqtPOMf
yNIrwL4mQUysbOZXC23SGH8rTrEgEFyQtN2m5aLrHd+9QLLY4t3IBB+227PIVcGuJLJThTOtPdew
xsS6yfXOUSW6apgWyDIfNjUrIg9L9dv8/WLneevnnsA5iOviaf+RUmO9TXQ/tkemP0H8isN13PoL
KRIVGQcqwBayLgVhXTKk2D4T/HxJFdkbNjrze7pMhgmXhDf+GbVyoRLOxGl5EDo1XBIw1mlL8d7m
xQXg0sQzbFhRd+KbXGiduXwLfLsrhq0hnyTT8HGwZiwoM4Kj9uNqTxoaLy289C332yX/mkmnm3mW
PD1qBz1oE0L9K5tlCfMERVbrQTORaV/BSimdkhaKlyXuwACIKJqBk4OX7jZbZ23oS2G2Wt5FHG0T
dtOcE9HrLiGMIVOpt19BjMKerMTy/wo22vcKE+I5TGlyiKRo/ZtZ3wK9sO+tmB1Zsyx4RGKa+kHp
4EzoC362MWXn1qjrtiqh0kFto6a0w1ftP/N6h6YEtDnUALkin6GJ/JoWpo++2xiWjqGxqEbd9ssf
DDLO/amL1sgWd8TlTI/NwktFggctxSk+6qzYgc0qH4EJkYWEI5XISyu9govWMBvqITdVU2d//B63
MkwFQ6Q64wInb20XI479okHFhXfjGTW1RuJmt63OowYFLFKrlVBYGYWJHKv9BMWo/ibMNtpcgUYx
SF++t+Up5KtbWJr/E5TClK3fGZP7QEgHG1Mf6m10UNJe1mQkTooNlktysXCFFD1YrIcmTzveDJ/k
xgIwSt+dNQWMZcwIeELcLfLRTpSQ0BwAqDifLd8DvE+VV8OlT3Z9juK9zYjzbqDBv7li3C6W9X6D
ExJl2WJPL8/N1RhaWg/1eHP8IL9NOxgE18APiNJ6Y9WUpJFsTqtx22wCQeQ3j0vduY35wU3pV8W8
g/P56qrK8AFy7GWBdw7ycadZuxXuyXbA0EISVgapyGLJVj/23NNBvopm0+/vhth3F2Wt8vU8zY5t
He0PhiRaY+YCD2oOgOERGTgl3AmYKmZUWu000RuYUEul7zsFOjn1+tWusHt0de0=
`protect end_protected
